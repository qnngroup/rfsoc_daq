`default_nettype none
`timescale 1ns / 1ps

module pwl_tb #(parameter SAMPLE_WIDTH, parameter DMA_DATA_WIDTH, parameter BATCH_SIZE)
					   (input wire clk,
					   	input wire valid_batch, 
					   	input wire[BATCH_SIZE-1:0][SAMPLE_WIDTH-1:0] batch,
					   	input wire pwl_rdy,
					   	output logic rst, 
					   	output logic halt, run_pwl,
					    Axis_IF dma);
	int period_len; 
	int expc_wave [$];
	logic clk2;
	assign clk2 = clk; 
	task automatic init();
		{halt, run_pwl} <= 0;
		{dma.data,dma.valid,dma.last} <= 0;
		sim_util_pkg::flash_signal(rst,clk2);
	endtask 

	function void clear_wave();
		while (expc_wave.size() > 0) expc_wave.pop_back();
		period_len = 0;
	endfunction

	function void reverse_wave();
		int expc_wave_tmp [$];
		while (expc_wave.size() > 0) expc_wave_tmp.push_back(expc_wave.pop_back());
	    expc_wave = expc_wave_tmp;
	endfunction

	task automatic halt_pwl();
		run_pwl <= 0;
		sim_util_pkg::flash_signal(halt,clk2);
	endtask

	task automatic send_buff(input logic[DMA_DATA_WIDTH-1:0] dma_buff [$], input bit osc_valid = 0, input int osc_delay_range[1:0] = {0,5});
		int delay_timer; 
		halt_pwl();
		while (~pwl_rdy) @(posedge clk); 
		for (int i = 0; i < dma_buff.size(); i++) begin
			dma.valid <= 1; 
			dma.data <= dma_buff[i]; 
			if (i == dma_buff.size()-1) dma.last <= 1; 
			@(posedge clk); 
			while (~dma.ready) @(posedge clk); 
			if (osc_valid) begin 
				{dma.valid,dma.last} <= 0; 
				@(posedge clk);
				delay_timer = $urandom_range(osc_delay_range[0],osc_delay_range[1]);
				repeat(delay_timer) @(posedge clk);				
			end 
		end
		{dma.valid,dma.last} <= 0; 
		@(posedge clk);		
	endtask 

	task automatic send_single_batch(input bit is_sparse, input bit is_fract, input bit is_neg); 
		logic[DMA_DATA_WIDTH-1:0] dma_buff [$];
		clear_wave();
		if (is_sparse) begin
			case ({is_fract,is_neg})
				2'b00: begin
					dma_buff = {64'd8589934625};
					expc_wave = {30,28,26,24,22,20,18,16,14,12,10,8,6,4,2,0};
				end 
				2'b01: begin
					dma_buff = {64'd35465799820902433};
					expc_wave = {-40,-29,-18,-7,4,15,26,37,48,59,70,81,92,103,114,125};
				end 
				2'b10: begin
					dma_buff = {64'd5840764961};
					expc_wave = {20,19,18,16,15,14,12,11,10,8,7,5,4,3,1,0};
				end 
				2'b11: begin
					dma_buff = {64'd3377679135146017};
					expc_wave = {-61,-56,-51,-47,-42,-37,-32,-27,-23,-18,-13,-8,-3,1,6,11};
				end 				
			endcase
		end else begin 
			case ({is_fract,is_neg})
				2'b00: begin
					dma_buff = {64'd8589934608, 64'd4503850882957316, 64'd37717504071565320, 64'd4294967298, 64'd281474976710658};
					expc_wave = {1,0,33,67,100,133,75,16,14,12,10,8,6,4,2,0};
				end 
				2'b01: begin
					dma_buff = {64'd281448133165072, 64'd18432670437156716558, 64'd37436171902517250};
					expc_wave = {133,107,81,55,28,2,-24,-50,-44,-37,-31,-25,-19,-12,-6,0};
				end 
				2'b10: begin
					dma_buff = {64'd3097951857541136, 64'd908878200820465668, 64'd319191411335364616, 64'd1406928206954498, 64'd18418596576038486018};
					expc_wave = {-100,4,286,569,851,1133,2181,3228,2826,2424,2022,1620,1217,815,413,11};
				end 
				2'b11: begin
					dma_buff = {64'd85899345930, 64'd28147497671065608, 64'd28428543151046660, 64'd18418596576038486022, 64'd18418597005535215618, 64'd2};
					expc_wave = {0,-100,-100,-100,-100,0,100,100,100,100,100,80,60,40,20,0};
				end 				
			endcase
		end 
		send_buff(dma_buff);
		period_len = 1; 
	endtask 

	task automatic send_pwl_wave(input bit osc_valid, input int osc_delay_range[1:0], input bit long_wave);
		logic[DMA_DATA_WIDTH-1:0] dma_buff [$];
		clear_wave();
		if (long_wave) begin 
			dma_buff = {64'd281294997160001, 64'd18069567424937721876, 64'd17951628349657120780, 64'd17464113689994264606, 64'd16244767985191878658, 64'd16418719520799064097, 64'd755200016804479000, 64'd2842894897700012040, 64'd2222242574053015617, 64'd15704893958493437958, 64'd15239617750855319578, 64'd14866381931736989729, 64'd14407014769745199114, 64'd14262922267812954130, 64'd8938800360205123588, 64'd8876594390352068737, 64'd6883470080263913490, 64'd6603118543320449038, 64'd5256542254736670849, 64'd11391570847122128910, 64'd10044721139929120786, 64'd13065229115011170322, 64'd16086010848604454926, 64'd14895371697118380065, 64'd12173790147303047176, 64'd11493187519535513624, 64'd12492423686858342561, 64'd706784937006465038, 64'd1289716537991692306, 64'd224896701095280737, 64'd12992601644690636820, 64'd11809284203747475468, 64'd12421210803116441729, 64'd500182589466738716, 64'd1927818225008836612, 64'd1417785567209128001, 64'd11705699585811546209, 64'd10854237781261811736, 64'd10641163613516201992, 64'd11196513742566326401, 64'd1637342058495737864, 64'd2193247884373262360, 64'd16602233417168453644, 64'd14583223649140736018, 64'd17595000526463500290, 64'd17577549077907439681, 64'd17016006499369680920, 64'd16805462818789785608, 64'd16630948333229179041, 64'd13140658622017044494, 64'd12835258495441502226, 64'd12574331192030724257, 64'd10254132959004786698, 64'd10108611668543668246, 64'd10707027469030523041, 64'd15058349134000553990, 64'd15221603724946374682, 64'd15165590204580954273, 64'd14821627783040532482, 64'd14817405164110413854, 64'd14267121584641081364, 64'd13900078668065013772, 64'd13858138896535126020, 64'd13843792828412067868, 64'd3699434667760025612, 64'd7257719531592744964, 64'd10926864502073393168, 64'd14023370720867319836, 64'd995617511347060738, 64'd3651292991395856386, 64'd3624552868608344225, 64'd1493224344955256850, 64'd1253688575746703374, 64'd808395162590445729, 64'd14166916082301468682, 64'd13848570064282845206, 64'd14720861017109168289, 64'd2618562918457802756, 64'd2777315295438438428, 64'd4337249616368893954, 64'd4448992401676435486, 64'd3386987314547130465, 64'd18435765469405642780, 64'd17444691614516838404, 64'd17242592581238587457, 64'd14008445098833149966, 64'd13300822370574598162, 64'd15554592509096820769, 64'd1114644728863457290, 64'd2366641699048259606, 64'd2435040118388949121, 64'd2833045735457816586, 64'd2864288814227980310, 64'd2468816471949508673, 64'd1317865292179636226, 64'd1281835791432417310, 64'd50664243300007969, 64'd17184046075677638684, 64'd16034783451085537284, 64'd15832121467853864993, 64'd14209699702093643800, 64'd12992605645838745608, 64'd13568221973212037217, 64'd2029155302958694426, 64'd3900115261054320646, 64'd3503798493845717185, 64'd9265034606286864481, 64'd4259565095441268766, 64'd8460291364180525058, 64'd8328561075079938081, 64'd6220032024540413974, 64'd4770436083013386250, 64'd4173427657410085025, 64'd13065788714026926209, 64'd2043228626037637128, 64'd2507650356767359000, 64'd12924476294875316232, 64'd10247378926584463384, 64'd10974428791428087937, 64'd14851746595617374238, 64'd15760630952348155906, 64'd15929797413351260225, 64'd2896661566717755402, 64'd3742491956622589974, 64'd4222688266890969217, 64'd7017171835674361860, 64'd7104709887153668124};
			expc_wave = {25241,25241,25241,25241,25241,25241,25241,25241,25241,25241,25241,25241,25241,25241,25085,24930,24775,24620,24465,24310,24155,24000,23844,23689,23534,23379,23224,23069,22914,22758,22603,22448,22293,22138,21983,21828,21673,21517,21362,21207,21052,20897,20742,20587,20432,20276,20121,19966,19811,19656,19501,19346,19191,19035,18880,18725,18570,18415,18260,18105,17949,17794,17639,17484,17329,17174,17019,16864,16708,16553,16398,16243,16088,15933,15778,15623,15467,15312,15157,15002,14847,14692,14537,14382,14227,14072,13917,13761,13606,13451,13296,12695,12094,11493,10892,10291,9690,9089,8488,7887,7286,6685,6084,5483,4882,4281,3680,3079,2478,1876,1275,674,73,-528,-1129,-1730,-2331,-2932,-3533,-4134,-4735,-5336,-5937,-6538,-7139,-7740,-8341,-8942,-9543,-9759,-9974,-10189,-10404,-10620,-10835,-11050,-11265,-11481,-11696,-11911,-12126,-12342,-12557,-12772,-12987,-13202,-13417,-13632,-13848,-14063,-14278,-14493,-14709,-14924,-15139,-15354,-15570,-15785,-16000,-16215,-16431,-16646,-16861,-17076,-17292,-17507,-17722,-17937,-18153,-18368,-18583,-18798,-19014,-19229,-19444,-19659,-19875,-20090,-20305,-20520,-20735,-20951,-21166,-21381,-21596,-21812,-22027,-22242,-22457,-22673,-22888,-23103,-23318,-23534,-23749,-23964,-24179,-24395,-24610,-24825,-25040,-25256,-25471,-25686,-25901,-26117,-26332,-26547,-26762,-26978,-27193,-27408,-27623,-27839,-28054,-28269,-28484,-28700,-28915,-29130,-26752,-24375,-21997,-19620,-17243,-14866,-12488,-10111,-7734,-5356,-2979,-601,1776,4153,6531,8908,8495,8083,7671,7259,6847,6435,6023,5611,5199,4787,4375,3962,3550,3138,2726,2314,1902,1490,1077,665,253,-159,-571,-983,-1395,-1807,-2220,-2632,-3044,-3456,-3868,-4280,-4692,-5104,-5517,-5929,-6341,-6753,-7165,-7577,-7989,-8402,-8814,-9226,-9638,-10050,-10462,-10874,-11286,-11699,-12111,-12523,-12935,-13347,-13759,-14171,-14584,-14996,-15408,-15820,-16232,-16644,-17056,-17468,-17881,-18293,-18705,-19117,-18692,-18268,-17844,-17419,-16995,-16571,-16147,-15722,-15298,-14874,-14449,-14025,-13601,-13177,-12752,-12328,-11904,-11480,-11055,-10631,-10207,-9782,-9358,-8934,-8510,-8085,-7661,-7237,-6812,-6388,-5964,-5540,-5115,-4691,-4267,-3842,-3418,-2994,-2570,-2145,-1721,-1297,-872,-448,-24,400,825,1249,1673,2098,2522,2946,3370,3795,4219,4643,5068,5492,5916,6340,6765,7189,7613,8037,8462,8886,9310,9735,10159,10583,11007,11432,11856,12280,12705,13129,13553,13977,14402,14826,15250,15674,16098,16523,16947,17415,17883,18352,18820,19288,19756,20224,20692,21161,21629,22097,22565,23033,23502,23970,24438,24906,25374,25843,26311,26779,27247,27715,28183,28652,29120,29588,30056,29061,28066,27071,26076,25082,24087,23092,22097,21102,20107,19112,18118,17123,16128,15133,14138,13143,12149,11154,10159,9164,8169,7174,6179,5185,4190,3195,2200,1205,210,-785,-1779,-2774,-3769,-4764,-5759,-6754,-7749,-8743,-9738,-10733,-11728,-12723,-13718,-14713,-15707,-16702,-17697,-18692,-19687,-20682,-21677,-22671,-23666,-24661,-25656,-26651,-27646,-28641,-29635,-30630,-31625,-32620,-32150,-31681,-31211,-30742,-30272,-29803,-29334,-28864,-28395,-27925,-27456,-26986,-26517,-26047,-25578,-25109,-24639,-24170,-23700,-23231,-22761,-22292,-21822,-21353,-20884,-20414,-19945,-19475,-19006,-18536,-18067,-17597,-17128,-16659,-16189,-15720,-15250,-14781,-14311,-13842,-13372,-12903,-12434,-11964,-11495,-11025,-10556,-10086,-9617,-9147,-8678,-8209,-7739,-7270,-6800,-6331,-5861,-5392,-4922,-4453,-3984,-3514,-3045,-2575,-2106,-1636,-1167,-697,-228,241,711,1180,1650,2119,2589,3058,3528,3997,4466,4936,5405,5875,6344,6814,7283,7753,8222,8691,9161,9630,10100,10569,11039,11508,11978,12447,12916,13386,13855,13344,12833,12322,11810,11299,10788,10277,9765,9254,8743,8232,7720,7209,6697,6186,5675,5164,4652,4141,3630,3118,2607,2096,1585,1073,562,51,-460,-972,-1483,-1994,-2505,-3017,-3528,-4039,-4550,-5062,-5573,-6084,-6596,-7107,-7618,-8129,-8641,-9152,-9663,-10174,-10686,-11197,-11708,-12219,-12731,-13242,-13753,-14264,-14776,-15287,-15798,-16309,-16821,-17332,-17843,-18354,-18866,-19377,-19017,-18656,-18296,-17936,-17576,-17215,-16855,-16495,-16135,-15774,-15414,-15054,-14694,-14333,-13973,-13613,-13253,-12892,-12532,-12172,-11812,-11451,-11091,-10731,-10371,-10010,-9650,-9290,-8930,-8570,-8278,-7986,-7695,-7403,-7112,-6820,-6528,-6237,-5945,-5653,-5362,-5070,-4779,-4487,-4195,-3904,-3612,-3320,-3029,-2737,-2446,-2154,-1862,-1571,-1279,-987,-696,-404,-113,179,470,762,1054,1345,1637,1928,2220,2512,2803,3095,3387,3678,3970,4261,4553,4681,4809,4937,5065,5192,5320,5448,5576,5703,5831,5959,6087,6215,6342,6470,6598,6726,6853,6981,7109,7237,7365,7492,7620,7748,7876,8003,8131,8259,8387,8514,8642,8770,8897,9025,9153,9281,9408,9536,9664,9792,9919,10047,10175,10153,10131,10109,10087,10065,10043,10020,9998,9976,9954,9932,9910,9888,9866,9844,9822,9800,9777,9755,9733,9711,9689,9667,9645,9623,9601,9579,9557,9534,9512,9490,9468,9446,9424,9402,9380,9358,9336,9314,9292,9269,9247,9225,9203,9181,9159,9137,9115,9093,9071,9049,9026,9004,8982,8960,8938,8916,8894,8872,8850,8828,8806,8784,8761,8739,8717,8695,8673,8651,8629,8607,8585,8563,8541,8518,8496,8474,8452,8430,8408,7519,6629,5739,4850,3960,3070,2180,1291,401,-489,-1378,-2268,-3158,-4047,-4937,-5827,-6716,-7606,-8496,-9385,-10275,-11165,-12054,-12944,-13834,-14723,-15613,-16503,-17392,-18282,-17923,-17564,-17205,-16846,-16487,-16128,-15769,-15410,-15050,-14691,-14332,-13973,-13614,-13255,-12896,-12537,-12178,-11819,-11460,-11101,-10742,-10383,-10024,-9665,-9306,-8947,-8588,-8229,-7869,-7510,-7151,-6792,-6433,-6074,-5715,-5356,-4997,-4638,-4279,-3920,-3561,-3310,-3058,-2807,-2555,-2304,-2052,-1801,-1549,-1298,-1046,-795,-543,-292,-40,211,463,714,966,1217,1469,1720,1972,2223,2475,2726,2978,3229,3481,3732,3984,4235,4487,4738,4990,5241,5493,5744,5996,6247,6499,6750,7002,7253,7505,7756,8008,8259,8511,8762,9014,9265,9517,9768,10020,10271,10523,10774,11026,11277,11529,11780,12032,12284,12535,12787,13038,13290,13541,13793,14044,14296,14547,14799,15050,15302,15553,15805,15409,15013,14617,14222,13826,13430,13034,12638,12242,11846,11450,11055,10659,10263,9867,9585,9303,9021,8740,8458,8176,7894,7613,7331,7049,6767,6486,6204,5922,5640,5359,5077,4795,4513,4232,3950,3668,3386,3105,2823,2541,2259,1978,1696,1414,1132,851,569,287,5,-276,-558,-840,-1122,-1403,-1685,-1967,-2249,-2530,-2812,-3094,-3376,-3657,-3939,-4221,-4503,-4784,-5066,-5348,-5630,-5911,-6193,-6475,-6757,-7038,-7320,-7602,-7884,-8165,-8447,-8729,-9011,-9292,-9574,-9856,-10138,-10419,-10701,-10983,-11265,-11546,-11828,-12110,-12392,-12673,-12955,-13237,-13518,-13800,-14082,-14364,-14645,-14927,-15209,-15491,-15772,-16054,-16336,-16110,-15884,-15658,-15432,-15206,-14980,-14754,-14528,-14303,-14077,-13851,-13625,-13399,-13173,-12947,-12721,-12495,-12269,-12043,-11817,-11591,-11365,-11139,-10913,-10687,-10461,-10235,-10009,-9783,-9557,-9331,-9105,-8879,-8653,-8427,-8201,-7975,-7749,-7524,-7298,-7072,-6846,-6620,-6394,-6168,-5942,-5716,-5490,-5264,-5038,-4812,-4586,-4360,-4134,-3908,-3682,-3456,-3230,-3004,-2778,-2552,-2326,-2100,-1874,-1648,-1422,-1196,-970,-744,-519,-293,-67,159,385,611,837,1063,1289,1515,1741,1967,2193,2419,2645,2871,3097,3323,3549,3775,4001,4227,4453,4547,4641,4736,4831,4925,5020,5115,5209,5304,5399,5494,5588,5683,5778,5872,5967,6062,6156,6251,6346,6440,6535,6629,6724,6819,6913,7008,7103,7197,7292,7387,7481,7576,7671,7765,7860,7954,8049,8144,8238,8333,8428,8522,8617,8712,8806,8901,8996,9090,9185,9280,9374,9469,9563,9658,9753,9847,9942,10037,10131,10226,10321,10415,10510,10605,10699,10794,10888,10983,11078,11172,11267,11362,11456,11551,11646,11740,11835,11930,12024,12119,12213,12308,12403,12497,12592,12687,12781,12876,12971,3537,2162,787,-588,-1964,-3339,-4714,-6089,-7464,-8839,-10214,-11590,-12965,-14340,-15715,-17090,-18465,-19840,-21215,-22591,-23966,-25341,-26716,-466,25784,23677,21570,19464,17357,15250,13143,11036,8929,6822,4716,2609,502,-1605,-3712,-5819,-7926,-10032,-12139,-14246,-16353,-16328,-16303,-16278,-16253,-16229,-16204,-16179,-16154,-16023,-15893,-15763,-15632,-15502,-15371,-15241,-15111,-14980,-14850,-14720,-14590,-14459,-14329,-14199,-14068,-13938,-13808,-13677,-13547,-13416,-13286,-13156,-13025,-12895,-12880,-12865,-12850,-12834,-12819,-12804,-12788,-12773,-12758,-12743,-12727,-12712,-12697,-12682,-12666,-12651,-12636,-12620,-12605,-12590,-12575,-12559,-12544,-12529,-12513,-12498,-12483,-12468,-12452,-12437,-12422,-12407,-12391,-12376,-12361,-12345,-12330,-12315,-12300,-12284,-12269,-12254,-12239,-12223,-12208,-12193,-12177,-12162,-12147,-12132,-12116,-12101,-12086,-12070,-12055,-12040,-12025,-12009,-11994,-11979,-11964,-11948,-11933,-11918,-11902,-11887,-11872,-11857,-11841,-11826,-11811,-11795,-11780,-11765,-11750,-11734,-11719,-11704,-11689,-11673,-11658,-11642,-11627,-11612,-11596,-11581,-11566,-11551,-11535,-11520,-11505,-11490,-11474,-11459,-11652,-11845,-12038,-12232,-12425,-12618,-12811,-13004,-13198,-13391,-13584,-13777,-13971,-14164,-14357,-14550,-14744,-14937,-15130,-15323,-15516,-15710,-15903,-16096,-16289,-16483,-16676,-16869,-17062,-17256,-17449,-17642,-17835,-18029,-18222,-18415,-18608,-18801,-18995,-19188,-19381,-19574,-19768,-19961,-20154,-20347,-20541,-20734,-20927,-21120,-21314,-21507,-21700,-21893,-22086,-22280,-22473,-22666,-22859,-23053,-23246,-23439,-23632,-23826,-24019,-24212,-24405,-24598,-24792,-24985,-25178,-25371,-25565,-25758,-25951,-26144,-26338,-26531,-26724,-26917,-27111,-27304,-27497,-27691,-27884,-28077,-28270,-28464,-28657,-28850,-29043,-29237,-29430,-29623,-29519,-29416,-29313,-29210,-29107,-29004,-28901,-28798,-28695,-28592,-28489,-28386,-28283,-28180,-28077,-27974,-27871,-27768,-27665,-27562,-27459,-27356,-27253,-27150,-27047,-26944,-26840,-26737,-26634,-26531,-26428,-26325,-26222,-26119,-26016,-25913,-25810,-25707,-25604,-25501,-25398,-25295,-25192,-25089,-24986,-24883,-24780,-24677,-24574,-24470,-24367,-24264,-24161,-24058,-23955,-23852,-23749,-23646,-23543,-23440,-23337,-23234,-23131,-23028,-22925,-22822,-22719,-22616,-22513,-22410,-22307,-22204,-22101,-21997,-21894,-21791,-21688,-21585,-21482,-21379,-21276,-21173,-21070,-20967,-20864,-20761,-20658,-20555,-20452,-20349,-20246,-20143,-20040,-19937,-19782,-19627,-19472,-19317,-19162,-19007,-18852,-18697,-18542,-18387,-18232,-18077,-17922,-17767,-17612,-17457,-17302,-17147,-16992,-16837,-16682,-16527,-16372,-16217,-16062,-15907,-15752,-15597,-15442,-15287,-15132,-14977,-14822,-14667,-14512,-14357,-14202,-14047,-13892,-13737,-13582,-13427,-13272,-13117,-12962,-12807,-12652,-12497,-12342,-12187,-12032,-11877,-11722,-11567,-11412,-11257,-11102,-10947,-10792,-10637,-10482,-10327,-10172,-10017,-9862,-9707,-9552,-9397,-9242,-9087,-8932,-8777,-8622,-8467,-8312,-8157,-8002,-7847,-7692,-7537,-7382,-7227,-7072,-6917,-6762,-6607,-6452,-6297,-6142,-5987,-5832,-5770,-5707,-5645,-5583,-5520,-5458,-5396,-5333,-5271,-5209,-5146,-5084,-5021,-4959,-4897,-4834,-4772,-4710,-4647,-4585,-4523,-4460,-4398,-4336,-4273,-4211,-4149,-4086,-4024,-3962,-3899,-3837,-3775,-3712,-3650,-3588,-3525,-3463,-3401,-3338,-3276,-3214,-3151,-3089,-3027,-4216,-5405,-6593,-7782,-8971,-10160,-11348,-12537,-13726,-12531,-11336,-10140,-8945,-7749,-6554,-5358,-4163,-2967,-1772,-577,619,1814,3009,4205,5400,6596,7791,7297,6804,6310,5817,5324,4830,4337,3844,3350,2857,2364,1870,1377,884,390,-103,-597,-1090,-1583,-2077,-2570,-3063,-3557,-4050,-4543,-5037,-5530,-6024,-6517,-7010,-7504,-7997,-8490,-8984,-9477,-9970,-10464,-10957,-11451,-11944,-12437,-12931,-13424,-13917,-14411,-14904,-15397,-15891,-16384,-16877,-17371,-17864,-18358,-18851,-19344,-19838,-20331,-20824,-21318,-21811,-22304,-22798,-23291,-23785,-24278,-24771,-25265,-25758,-26251,-26744,-27238,-27731,-27668,-27605,-27542,-27479,-27416,-27353,-27290,-27227,-27164,-27101,-27038,-26975,-26912,-26849,-26786,-26723,-26660,-26597,-26534,-26471,-26408,-26345,-26282,-26219,-26156,-26093,-26030,-25967,-25904,-25840,-25777,-25714,-25651,-25588,-25525,-25462,-25399,-25336,-25273,-25210,-25147,-25084,-25021,-24958,-24895,-24832,-24769,-24706,-24643,-24580,-24517,-24454,-24391,-24328,-24265,-24202,-24139,-24076,-24013,-23950,-23045,-22139,-21233,-20327,-19421,-18515,-17610,-16704,-15798,-14892,-13986,-13080,-12175,-11269,-10363,-9457,-8551,-7646,-6740,-5834,-4928,-4022,-3116,-2211,-1305,-399,507,1413,2319,3224,4130,5036,5942,6848,6486,6124,5762,5400,5037,4675,4313,3951,3588,3226,2864,2502,2139,1777,1415,1053,690,328,-34,-396,-759,-1121,-1483,-1845,-2208,-2570,-2932,-3294,-3657,-4019,-4381,-4743,-5106,-5468,-5830,-6192,-6555,-6917,-7279,-7641,-8004,-8366,-8728,-9090,-9453,-9815,-10177,-10539,-10902,-11264,-11626,-11988,-12351,-12713,-13075,-13437,-13800,-14162,-14524,-14886,-15249,-15611,-15973,-16335,-16698,-17060,-17422,-17784,-18147,-18509,-18871,-19233,-19596,-19958,-20320,-20682,-21045,-21407,-21770,-22132,-22494,-22856,-23219,-23581,-23161,-22741,-22320,-21900,-21480,-21059,-20639,-20219,-19798,-19378,-18957,-18537,-18117,-17696,-17276,-16856,-16435,-16015,-15595,-15174,-14754,-14334,-13913,-13493,-13073,-12653,-12232,-11812,-11392,-10971,-10551,-10131,-9710,-9290,-8870,-8449,-8029,-7609,-7188,-6768,-6348,-5927,-5507,-5087,-4666,-4246,-3826,-3405,-2985,-2565,-2144,-1724,-1304,-883,-463,-43,378,798,1218,1639,2059,2479,2900,3320,3740,4161,4581,4286,3990,3694,3398,3103,2807,2511,2215,1919,1623,1327,1032,736,440,144,-152,-447,-743,-1039,-1335,-1631,-1926,-2222,-2518,-2814,-3110,-3406,-3701,-3997,-4293,-4589,-4885,-5180,-5476,-5772,-6068,-6364,-6659,-6955,-7251,-7547,-7843,-8138,-8434,-8730,-9026,-9322,-9617,-9913,-10209,-10505,-10801,-11097,-11392,-11688,-11984,-12280,-12576,-12871,-13167,-13463,-13759,-14055,-14350,-14646,-14942,-15238,-15534,-15829,-16125,-16421,-16717,-17013,-17308,-17604,-17900,-18196,-18492,-18788,-19083,-19379,-19675,-19971,-20267,-20562,-20858,-21154,-21450,-21746,-22042,-22338,-22633,-22929,-23225,-23521,-23817,-24112,-24408,-24704,-24100,-23496,-22891,-22287,-21682,-21078,-20474,-19870,-19265,-18661,-18057,-17452,-16848,-16244,-15639,-15035,-14431,-13827,-13222,-12618,-12014,-11409,-10805,-10201,-9597,-8992,-8388,-9580,-10773,-11965,-13157,-14350,-15542,-16734,-17927,-19119,-20311,-21504,-22696,-23888,-25081,-26273,-27465,-28658,-29850,-29167,-28483,-27800,-27116,-26433,-25749,-25066,-24382,-23699,-23016,-22332,-21649,-20965,-20282,-19598,-18915,-18232,-17548,-16865,-16181,-15498,-14814,-14131,-13447,-12764,-12081,-11397,-10714,-10030,-9347,-8663,-7980,-7297,-6613,-5930,-5246,-4563,-3879,-3196,-2513,-1829,-1146,-462,221,905,1588,2272,2955,3638,4322,5005,5689,6372,7056,7739,8422,9106,9789,10473,11156,11840,12523,13207,13890,14573,15257,15940,16624,17307,17991,18674,19357,20041,20724,21408,22091,22775,23458,23569,23680,23790,23901,24011,24122,24233,24343,24454,24565,24675,24786,24897,25007,25118,25229,25339,25450,25560,25671,25782,25892,26003,26114,26224,26335,26446,26556,26667,26777,26888,26999,27109,27220,27331,27441,27552,27663,27773,27884,27995,28105,28216,28326,28437,28548,28658,28769,28880,28990,29101,29212,29322,29433,29543,29654,29765,29875,29986,30097,30207,30318,30429,30539,30650,30761,30871,30982,31092,31203,31314,31424,31535,31645,31756,26576,21396,16216,11036,5856,676,-4504,-9684,-14864,-14761,-14659,-14557,-14455,-14353,-14251,-14149,-14047,-13945,-13843,-13741,-13639,-13537,-13435,-13333,-13231,-13129,-13027,-12925,-12823,-12721,-12619,-12517,-12415,-12313,-12211,-12109,-12007,-11905,-11803,-11701,-11599,-11497,-11395,-10844,-10293,-9742,-9191,-8640,-8089,-7538,-6986,-6435,-5884,-5333,-4782,-4231,-3680,-3129,-2577,-2026,-1475,-924,-373,178,729,1280,1832,2383,2934,3485,4036,4587,5138,5689,6241,6792,7343,7894,8446,8997,9548,10099,9481,8863,8245,7627,7009,6391,5773,5155,4537,3919,3301,2683,2065,1447,829,211,-407,-1025,-1643,-2261,-2879,-3497,-4115,-4733,-5351,-5969,-6587,-7205,-7823,-7534,-7245,-6957,-6668,-6379,-6090,-5802,-5513,-5224,-4936,-4647,-4358,-4069,-3781,-3492,-3204,-2915,-2626,-2337,-2049,-1760,-1718,-1676,-1634,-1592,-1551,-1509,-1467,-1425,-1383,-1341,-1299,-1257,-1215,-1173,-1131,-1090,-1048,-1006,-964,-922,-880,-838,-796,-754,-712,-670,-629,-587,-545,-503,-461,-419,-377,-335,-293,-251,-210,-168,-126,-84,-42,0};
		end else begin 
			dma_buff = {64'd281469822763018, 64'd18445055228534718486, 64'd1688850576113697, 64'd2533275506245648, 64'd3096222954225680, 64'd2251798024093729, 64'd4294967316, 64'd3096214006398988, 64'd18445618163065290760, 64'd18442521951393087512, 64'd18444492276230062145, 64'd2533277124591620, 64'd3096216153882634, 64'd18};
			expc_wave = {0,0,0,0,0,0,0,0,0,2,4,6,8,10,10,9,9,8,8,7,7,6,6,5,4,4,3,3,2,2,1,1,0,0,-1,-1,-2,-3,-3,-4,-4,-5,-5,-6,-6,-7,-7,-8,-9,-10,-10,-11,-11,-12,-12,-13,-13,-14,-14,-15,-12,-10,-7,-5,-2,0,3,5,8,10,9,8,7,6,5,4,3,2,1,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,7,7,7,8,8,9,9,10,10,10,10,10,10,10,9,9,9,9,8,8,8,8,8,8,7,7,7,7,7,7,6,6,6,5,4,3,2,1,-1,-2,-3,-4,-5,-6,-5,-4,-2,-1,0};
		end 
		send_buff(dma_buff, osc_valid, osc_delay_range);
		period_len = expc_wave.size()/BATCH_SIZE;
	endtask  					   

	task automatic check_pwl_wave(inout sim_util_pkg::debug debug, input int periods_to_check);
		int expc_wave_tmp [$];
		int samples_seen,periods_seen,expc_sample;
		bit do_print;
		string err_str;
		periods_seen = 0; 
		run_pwl <= 1; 
		@(posedge clk);
		repeat(periods_to_check) begin
			expc_wave_tmp = expc_wave;
			samples_seen = 0; 
			debug.displayc($sformatf("\nPeriod %0d",periods_seen), .msg_color(sim_util_pkg::BLUE), .msg_verbosity(sim_util_pkg::DEBUG));
			for (int i = 0; i < period_len; i++) begin
				while (~valid_batch) @(posedge clk); 
				for (int j = 0; j < BATCH_SIZE; j++) begin 
					expc_sample = expc_wave_tmp.pop_back();
					if (expc_wave.size() > 300) begin
						if ($signed(batch[j]) != expc_sample) do_print = 1; 
						else if (j == 15) do_print = 1;
						else do_print = 0;
						err_str = (debug.get_error_count() > 100)? "." : $sformatf("Error on %0dth sample: Expected %0d, Got %0d",samples_seen, expc_sample, $signed(batch[j]));
						if (do_print) debug.disp_test_part(1+samples_seen, $signed(batch[j]) == expc_sample,err_str);
					end else debug.disp_test_part(1+samples_seen, $signed(batch[j]) == expc_sample,$sformatf("Error on %0dth sample: Expected %0d, Got %0d",samples_seen, expc_sample, $signed(batch[j])));
					samples_seen++;
				end 
				@(posedge clk); 
			end
			periods_seen++;
		end
	endtask 
endmodule 

`default_nettype wire

