// Axis_If.sv - Reed Foster
// single axi-stream interface
interface Axis_If #(
  parameter DWIDTH = 32
);

logic [DWIDTH - 1:0]  data;
logic                 ready;
logic                 valid;
logic                 last;
logic                 ok;

assign ok = ready & valid;

// master/slave packetized interface
modport Master (
  input   ready,
  output  valid,
  output  data,
  output  last,
  input   ok
);

modport Slave (
  output  ready,
  input   valid,
  input   data,
  input   last,
  input   ok
);

/* verilator lint_off MULTIDRIVEN */

////////////////////////////////
// Utitlities for testbenches //
////////////////////////////////

// Combined with a process that updates data_in whenever
// ok = valid && ready is high, this task sends samples to
// an Axis_If interface.
// Can optionally toggle the valid signal randomly to test
// handshaking logic of modules
task automatic send_samples(
  ref clk, // reference to clock signal in testbench
  input int n_samples, // number of samples to send
  input bit rand_arrivals, // if 1, toggle valid, otherwise leave it high
  input bit reset_valid // if 1, reset valid signal after sending the samples
);
  int samples_sent;
  // reset
  samples_sent = 0;
  valid <= 1'b1;
  while (samples_sent < n_samples) begin
    @(posedge clk);
    if (ok) begin
      samples_sent = samples_sent + 1'b1;
    end
    if (rand_arrivals) begin
      valid <= 1'($urandom()) & 1'b1;
    end // else do nothing; intf.valid is already 1'b1
  end
  if (reset_valid) begin
    valid <= '0;
    @(posedge clk);
  end
endtask

// Update registers with an Axis_If interface
// must be augmented with a process or other statement to actually update the
// data
task automatic send_sample_with_timeout(
  ref clk,
  input int timeout,
  output logic success
);
  int timer;
  timer = 0;
  success = 1'b0;
  valid <= 1'b1;
  while ((timer < timeout) & (~success)) begin
    timer = timer + 1;
    if (ok) begin
      success = 1'b1;
    end
    @(posedge clk);
  end
  valid <= 1'b0;
endtask


// Wait until the last transfer goes through on an Axis_If interface,
// or until a timeout is reached. Can optionally toggle the ready signal
// to test backpressure handling logic of modules
task automatic do_readout(
  ref clk, // reference to clock signal in testbench
  input bit rand_ready, // if 1, toggle ready, otherwise leave it high
  input int timeout // number of clock cycles to wait for if last is never asserted
);
  int cycle_count;
  cycle_count = 0;
  ready <= 1'b0;
  // wait a bit before actually doing the readout
  repeat (500) @(posedge clk);
  ready <= 1'b1;
  // give up after timeout clock cycles if last is not achieved
  while ((!(last & ok)) & (cycle_count < timeout)) begin
    @(posedge clk);
    cycle_count = cycle_count + 1;
    if (rand_ready) begin
      ready <= 1'($urandom()) & 1'b1;
    end
  end
  @(posedge clk);
  ready <= 1'b0;
endtask

/* verilator lint_on MULTIDRIVEN */

endinterface
