// sparse_sample_buffer_test.sv - Reed Foster
// Check that the combined banked sample_buffer and sample_discriminator work
// correctly, saving the correct data and outputting it in the correct format
// (i.e. timestamps first, then data, and for each bank, outputting the
// corresponding channel index and sample quantity stored in that bank)

`timescale 1ns / 1ps
module sparse_sample_buffer_test ();

sim_util_pkg::math #(int) math; // abs, max functions on integers
sim_util_pkg::debug debug = new(sim_util_pkg::DEFAULT); // printing, error tracking

logic clk = 0;
localparam CLK_RATE_HZ = 100_000_000;
always #(0.5s/CLK_RATE_HZ) clk = ~clk;

logic reset;

localparam int CHANNELS = 8;
localparam int TSTAMP_BUFFER_DEPTH = 128;
localparam int DATA_BUFFER_DEPTH = 1024;
localparam int AXI_MM_WIDTH = 128;
localparam int PARALLEL_SAMPLES = 4;
localparam int SAMPLE_WIDTH = 16;
localparam int APPROX_CLOCK_WIDTH = 48;

// derived parameters
localparam int SAMPLE_INDEX_WIDTH = $clog2(DATA_BUFFER_DEPTH*CHANNELS);
localparam int TIMESTAMP_WIDTH = SAMPLE_WIDTH * ((SAMPLE_INDEX_WIDTH + APPROX_CLOCK_WIDTH + (SAMPLE_WIDTH - 1)) / SAMPLE_WIDTH);

// util for parsing timestamp/sample data from buffer output
sparse_sample_buffer_pkg::util #(
  .AXI_MM_WIDTH(AXI_MM_WIDTH),
  .TIMESTAMP_WIDTH(TIMESTAMP_WIDTH),
  .SAMPLE_WIDTH(SAMPLE_WIDTH),
  .PARALLEL_SAMPLES(PARALLEL_SAMPLES),
  .DATA_BUFFER_DEPTH(DATA_BUFFER_DEPTH),
  .CHANNELS(CHANNELS)
) buf_util;

Realtime_Parallel_If #(.DWIDTH(PARALLEL_SAMPLES*SAMPLE_WIDTH), .CHANNELS(CHANNELS)) data_in ();
Axis_If #(.DWIDTH(AXI_MM_WIDTH)) data_out ();
Axis_If #(.DWIDTH($clog2($clog2(CHANNELS)+1))) buffer_config ();
Axis_If #(.DWIDTH(2)) buffer_start_stop ();
Axis_If #(.DWIDTH(CHANNELS*SAMPLE_WIDTH*2)) sample_discriminator_config();

logic capture_start, capture_stop, start_aux;
logic [$clog2($clog2(CHANNELS)+1)-1:0] banking_mode;
logic [CHANNELS-1:0][SAMPLE_WIDTH-1:0] threshold_high, threshold_low;
logic capture_done;

always_comb begin
  for (int i = 0; i < CHANNELS; i++) begin
    sample_discriminator_config.data[2*SAMPLE_WIDTH*i+:2*SAMPLE_WIDTH] = {threshold_high[i], threshold_low[i]};
  end
end

assign buffer_config.data = banking_mode;
assign buffer_start_stop.data = {capture_start, capture_stop};

sparse_sample_buffer #(
  .CHANNELS(CHANNELS),
  .TSTAMP_BUFFER_DEPTH(TSTAMP_BUFFER_DEPTH),
  .DATA_BUFFER_DEPTH(DATA_BUFFER_DEPTH),
  .AXI_MM_WIDTH(AXI_MM_WIDTH),
  .PARALLEL_SAMPLES(PARALLEL_SAMPLES),
  .SAMPLE_WIDTH(SAMPLE_WIDTH),
  .APPROX_CLOCK_WIDTH(APPROX_CLOCK_WIDTH)
) dut_i (
  .clk,
  .reset,
  .timestamp_width(),
  .capture_done,
  .data_in,
  .data_out,
  .sample_discriminator_config,
  .buffer_config,
  .buffer_start_stop,
  .start_aux
);

// allow the data to be manually updated when we change the range so the first sample for a new range isn't stale
// this simplifies the testing
logic update_input_data;
logic [CHANNELS-1:0][SAMPLE_WIDTH-1:0] data_range_low, data_range_high;
logic [PARALLEL_SAMPLES*SAMPLE_WIDTH-1:0] data_sent [CHANNELS][$];
logic [AXI_MM_WIDTH-1:0] data_received [$];
int last_received [$];
logic [CHANNELS-1:0][TIMESTAMP_WIDTH-SAMPLE_INDEX_WIDTH-1:0] timer;

// send data to DUT and save sent/received data
always @(posedge clk) begin
  for (int channel = 0; channel < CHANNELS; channel++) begin
    if (reset) begin
      data_in.data[channel] <= '0;
    end else begin
      if (data_in.valid[channel]) begin
        // save data that was sent
        data_sent[channel].push_front(data_in.data[channel]);
      end
      if (data_in.valid[channel] || update_input_data) begin
        // send new data
        for (int sample = 0; sample < PARALLEL_SAMPLES; sample++) begin
          data_in.data[channel][sample*SAMPLE_WIDTH+:SAMPLE_WIDTH] <= $urandom_range(data_range_low[channel], data_range_high[channel]);
        end
      end
    end
  end
  // save all data in the same buffer and postprocess it later
  if (data_out.ok) begin
    data_received.push_front(data_out.data);
    if (data_out.last) begin
      last_received.push_front(data_received.size());
    end
  end
end

task check_results(
  input int banking_mode,
  input logic [CHANNELS-1:0][SAMPLE_WIDTH-1:0] threshold_high,
  input logic [CHANNELS-1:0][SAMPLE_WIDTH-1:0] threshold_low,
  inout logic [CHANNELS-1:0][TIMESTAMP_WIDTH-SAMPLE_INDEX_WIDTH-1:0] timer,
  input int max_transfer_count,
  input bit buffer_filled
);
  // checks that:
  // - timestamps line up with when samples were sent
  // - all inputs > threshold_high were saved and all inputs < threshold_low
  //    were not
  // - all samples < threshold_high that were saved arrived in sequence after
  //    a sample > threshold_high

  // data structures for organizing DMA output
  logic [TIMESTAMP_WIDTH-1:0] timestamps [CHANNELS][$];
  logic [SAMPLE_WIDTH*PARALLEL_SAMPLES-1:0] samples [CHANNELS][$];

  // first report the size of the buffers
  for (int i = 0; i < CHANNELS; i++) begin
    debug.display($sformatf("data_sent[%0d].size() = %0d", i, data_sent[i].size()), sim_util_pkg::VERBOSE);
  end
  debug.display($sformatf("data_received.size() = %0d", data_received.size()), sim_util_pkg::VERBOSE);

  // make sure that last arrived before max_transfer_count samples
  if (last_received.size() !== 1) begin
    debug.error($sformatf(
      "expected a single tlast event, got %0d",
      last_received.size())
    );
  end else begin
    if (last_received[$] > max_transfer_count) begin
      debug.error($sformatf(
        "expected tlast event after at most %0d transfers, got it on the %0d transfer",
        max_transfer_count,
        last_received[$])
      );
    end
  end
  while (last_received.size() > 0) last_received.pop_back();

  ///////////////////////////////////////////////////////////////////
  // organize DMA output into data structures for easier analysis
  ///////////////////////////////////////////////////////////////////
  buf_util.parse_buffer_output(data_received, timestamps, samples);
  debug.display("parsed data_received:", sim_util_pkg::VERBOSE);
  for (int i = 0; i < CHANNELS; i++) begin
    debug.display($sformatf("timestamps[%0d].size() = %0d", i, timestamps[i].size()), sim_util_pkg::VERBOSE);
    debug.display($sformatf("samples[%0d].size() = %0d", i, samples[i].size()), sim_util_pkg::VERBOSE);
  end

  //////////////////////////////////////
  // process data "like normal"
  //////////////////////////////////////
  buf_util.check_timestamps_and_data(
    debug,
    banking_mode,
    threshold_high,
    threshold_low,
    timer,
    timestamps,
    samples,
    data_sent,
    buffer_filled
  );

endtask

task set_banking_mode(input int mode);
  banking_mode <= mode;
  buffer_config.valid <= 1'b1;
  while (~buffer_config.ok) @(posedge clk);
  buffer_config.valid <= 1'b0;
endtask

task start_acq(input bit use_axis);
  if (use_axis) begin
    capture_stop <= 1'b0;
    capture_start <= 1'b1;
    buffer_start_stop.valid <= 1'b1;
    @(posedge clk);
    capture_start <= 1'b0;
    buffer_start_stop.valid <= 1'b0;
  end else begin
    start_aux <= 1'b1;
    @(posedge clk);
    start_aux <= 1'b0;
  end
endtask

task stop_acq();
  capture_stop <= 1'b1;
  capture_start <= 1'b0;
  buffer_start_stop.valid <= 1'b1;
  @(posedge clk);
  capture_stop <= 1'b0;
  buffer_start_stop.valid <= 1'b0;
endtask

int samples_to_send;

initial begin
  debug.display("### RUNNING TEST FOR SPARSE_SAMPLE_BUFFER ###", sim_util_pkg::DEFAULT);
  reset <= 1'b1;
  capture_start <= 1'b0;
  capture_stop <= 1'b0;
  start_aux <= '0;
  timer <= '0; // reset timer for all channels
  banking_mode <= '0; // only enable channel 0 to start
  data_out.ready <= '0;
  data_in.valid <= '0;
  buffer_config.valid <= 1'b0;
  sample_discriminator_config.valid <= 1'b0;
  buffer_start_stop.valid <= 1'b0;
  repeat (100) @(posedge clk);
  reset <= 1'b0;
  repeat (50) @(posedge clk);
  
  for (int start_type = 0; start_type < 2; start_type++) begin
    for (int in_valid_rand = 0; in_valid_rand < 2; in_valid_rand++) begin
      for (int bank_mode = 0; bank_mode < 4; bank_mode++) begin
        set_banking_mode(bank_mode);
        for (int amplitude_mode = 0; amplitude_mode < 5; amplitude_mode++) begin
          repeat (10) @(posedge clk);
          unique case (amplitude_mode)
            0: begin
              // save everything
              for (int i = 0; i < CHANNELS; i++) begin
                data_range_low[i] <= 16'h03c0;
                data_range_high[i] <= 16'h04ff;
                threshold_low[i] <= 16'h0000;
                threshold_high[i] <= 16'h0100;
              end
            end
            1: begin
              // send stuff straddling the threshold with strong hysteresis
              for (int i = 0; i < CHANNELS; i++) begin
                data_range_low[i] <= 16'h00ff;
                data_range_high[i] <= 16'h04ff;
                threshold_low[i] <= 16'h01c0;
                threshold_high[i] <= 16'h0400;
              end
            end
            2: begin
              // send stuff below the threshold
              for (int i = 0; i < CHANNELS; i++) begin
                data_range_low[i] <= 16'h0000;
                data_range_high[i] <= 16'h01ff;
                threshold_low[i] <= 16'h0200;
                threshold_high[i] <= 16'h0200;
              end
            end
            3: begin
              // send stuff straddling the threshold with weak hysteresis
              for (int i = 0; i < CHANNELS; i++) begin
                data_range_low[i] <= 16'h0000;
                data_range_high[i] <= 16'h04ff;
                threshold_low[i] <= 16'h03c0;
                threshold_high[i] <= 16'h0400;
              end
            end
            4: begin
              // send stuff that mostly gets filtered out
              for (int i = 0; i < CHANNELS; i++) begin
                data_range_low[i] <= 16'h0000;
                data_range_high[i] <= 16'h04ff;
                threshold_low[i] <= 16'h03c0;
                threshold_high[i] <= 16'h0400;
              end
            end
          endcase
          // write the new threshold to the discriminator and update the input data
          sample_discriminator_config.valid <= 1'b1;
          update_input_data <= 1'b1;
          @(posedge clk);
          sample_discriminator_config.valid <= 1'b0;
          update_input_data <= 1'b0;

          repeat (10) @(posedge clk);
          start_acq(start_type & 1'b1);

          if (amplitude_mode == 0) begin
            // send enough samples to fill up buffer exactly
            samples_to_send = DATA_BUFFER_DEPTH*(8 >> bank_mode);
          end else begin
            samples_to_send = $urandom_range(50,500);
          end

          data_in.send_samples(clk, samples_to_send - 10, in_valid_rand & 1'b1, 1'b1);
          if (start_type === 1'b0) begin
            // retrigger start to make sure we can't accidentally trigger over
            // the current capture before it's read out
            start_acq(1'b0);
          end
          data_in.send_samples(clk, 10, in_valid_rand & 1'b1, 1'b1);
          repeat (10) @(posedge clk);
          if (amplitude_mode == 0) begin
            // check that capture_done is asserted
            if (capture_done !== 1'b1) begin
              debug.error("expected capture to be done, but it's not");
              stop_acq();
            end
          end else begin
            stop_acq();
          end
          repeat (10) @(posedge clk);
          if (start_type === 1'b0) begin
            // retrigger start to make sure we can't accidentally retrigger
            // capture before readout of the previous capture
            start_acq(1'b0);
          end
          repeat (10) @(posedge clk);
          data_out.do_readout(clk, 1'b1, 100000);
          debug.display($sformatf("checking results amplitude_mode = %0d", amplitude_mode), sim_util_pkg::VERBOSE);
          debug.display($sformatf("banking mode                    = %0d", bank_mode), sim_util_pkg::VERBOSE);
          debug.display($sformatf("samples sent with rand_valid    = %0d", in_valid_rand), sim_util_pkg::VERBOSE);
          check_results(
            bank_mode,
            threshold_high,
            threshold_low,
            timer,
            samples_to_send*(1 << bank_mode) + 2*CHANNELS + TSTAMP_BUFFER_DEPTH*(1 << bank_mode) + 2*CHANNELS,
            amplitude_mode == 0 
          );
        end
      end
    end
  end
  debug.finish();
end

endmodule
