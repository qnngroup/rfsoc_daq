`default_nettype none
`timescale 1ns / 1ps



module integrated_tb #(parameter BUS_WIDTH, parameter DATA_WIDTH)
					   (input wire clk, rst,
					    Recieve_Transmit_IF intf);
	

endmodule 

`default_nettype wire

