// axis_x2.sv - Reed Foster
// computes x^2 on axi-stream data
module axis_x2 #(
  parameter int SAMPLE_WIDTH = 16,
  parameter int PARALLEL_SAMPLES = 1,
  parameter int SAMPLE_FRAC_BITS = 16
) (
  input wire clk, reset,
  Axis_If.Slave data_in,
  Axis_If.Master data_out
);

// register signals to infer DSP hardware multiplier
// lots of pipeline registers to enable the DSP to run at high clock rates
// can't do packed arrays because of signed type
logic signed [SAMPLE_WIDTH-1:0] data_in_reg [PARALLEL_SAMPLES]; // 0Q16, 2Q14
// register the full-width product
logic signed [2*SAMPLE_WIDTH-1:0] product [PARALLEL_SAMPLES]; // 0Q32, 4Q28
// shift and truncate the product and register it
logic signed [SAMPLE_WIDTH-1:0] product_d [PARALLEL_SAMPLES]; // 0Q16, 4Q12
logic [3:0] valid_d, last_d;

always_ff @(posedge clk) begin
  if (reset) begin
    valid_d <= '0;
  end else begin
    if (data_in.ok) begin
      for (int i = 0; i < PARALLEL_SAMPLES; i++) begin
        data_in_reg[i] <= data_in.data[i*SAMPLE_WIDTH+:SAMPLE_WIDTH]; // 0Q16, 2Q14
      end
    end
    if (data_out.ready || (!data_out.valid)) begin
      for (int i = 0; i < PARALLEL_SAMPLES; i++) begin
        product[i] <= data_in_reg[i]*data_in_reg[i]; // 0Q16*0Q16 = 0Q32, 2Q14*2Q14 = 4Q28
        product_d[i] <= product[i][2*SAMPLE_WIDTH-1-:SAMPLE_WIDTH]; // 0Q16, 4Q12
        data_out.data[i*SAMPLE_WIDTH+:SAMPLE_WIDTH] <= product_d[i];
      end
      valid_d <= {valid_d[2:0], data_in.ok};
      last_d <= {last_d[2:0], data_in.last};
    end
  end
end

assign data_out.valid = valid_d[3];
assign data_out.last = last_d[3];
assign data_in.ready = data_out.ready;

endmodule
