// receive_top_test.sv - Reed Foster
// verifies data from ADC is saved correctly

