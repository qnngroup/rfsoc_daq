// awg_test.sv - Reed Foster

`timescale 1ns/1ps;

module awg_test ();
endmodule
