`default_nettype none
`timescale 1ns / 1ps
import mem_layout_pkg::*;

module top_level_tb #(parameter VERBOSE = 1)(input wire start, output logic[1:0] done);
    localparam TOTAL_TESTS = 3; 
    localparam STARTING_TEST = 0; 
    localparam TIMEOUT = 10_000; 
    localparam PERIODS_TO_CHECK = 3; 
    logic clk, rst;
    logic[15:0] timer; 

    enum logic[2:0] {IDLE, TEST, WRESP, CHECK, DONE} testState; 
    logic[1:0] test_check; // test_check[0] = check, test_check[1] == 1 => test passed else test failed 
    logic[7:0] test_num; 
    logic[7:0] testsPassed, testsFailed; 
    logic kill_tb; 
    logic panic = 0; 

    logic[`A_BUS_WIDTH-1:0] raddr_packet, waddr_packet;
    logic[`WD_BUS_WIDTH-1:0] rdata_packet, wdata_packet;
    logic[`DMA_DATA_WIDTH-1:0] pwl_tdata;
    logic[3:0] pwl_tkeep;
    logic pwl_tlast, pwl_tready, pwl_tvalid; 
    logic raddr_valid_packet, waddr_valid_packet, wdata_valid_packet, rdata_valid_out, wresp_valid_out, rresp_valid_out;
    logic ps_wresp_rdy,ps_read_rdy; 
    logic[1:0] wresp_out, rresp_out; 
    logic[(`BATCH_WIDTH)-1:0] dac_batch;
    logic valid_dac_batch, dac0_rdy;
    logic pl_rstn;
    logic[`BATCH_SAMPLES-1:0][`SAMPLE_WIDTH-1:0] init_samples, dac_samples;

    enum logic[1:0] {IDLE_PWL, SEND_BUFF,VERIFY} pwlTestState; 
    logic[$clog2(BUFF_LEN):0] dma_i;
    logic[$clog2(`PWL_BRAM_DEPTH):0] exp_i;
    logic send_dma_buff,run_pwl; 
    logic checked_full_wave;
    logic[$clog2(PERIODS_TO_CHECK):0] periods; 
    logic[`BATCH_SAMPLES-1:0][`SAMPLE_WIDTH-1:0] curr_expected_batch;
    logic[`BATCH_SAMPLES-1:0] error_vec;

    //DMA BUFFER TO SEND
    localparam BUFF_LEN = 67;
    logic[BUFF_LEN-1:0][`DMA_DATA_WIDTH-1:0] dma_buff;
    assign dma_buff = {48'h3c34097f0000, 48'h3b282a75ffe1, 48'h3a182a8dffff, 48'h390604140024, 48'h375602700001, 48'h36cb3a3eff99, 48'h36703d79fff7, 48'h34f71d030016, 48'h3443346affdf, 48'h327104f3001a, 48'h324d040c0006, 48'h31131b68ffed, 48'h31120d650e03, 48'h301c1123fffc, 48'h2f260edc0002, 48'h2cfb1f57fff8, 48'h2c6c0674002d, 48'h2c6b2764df10, 48'h2ba30ca90022, 48'h2ad63ceaffc4, 48'h28b9275b000a, 48'h288e1e7f0035, 48'h279d0edb0011, 48'h26383550ffe4, 48'h263737bcfd94, 48'h24212bb10006, 48'h238622e0000f, 48'h23762622ffcc, 48'h220302a70018, 48'h21d22479ff4f, 48'h203a0b6d0010, 48'h1f670a900001, 48'h1e4b29f8ffe4, 48'h1e4a07bb223d, 48'h1d023937ffd9, 48'h1c2328e40013, 48'h1b1337a5fff2, 48'h1aab3907fffd, 48'h1a0c353f0006, 48'h18843a7efffd, 48'h17451c9c0018, 48'h171d2593ffc7, 48'h161e2d7ffff8, 48'h13cd06900011, 48'h12de066d0001, 48'h126c10d1ffe9, 48'h11732742ffe9, 48'h11720a321d10, 48'h105a01ec0008, 48'hfc72405ffc5, 48'he801dfd0005, 48'hd2a18a40004, 48'hc1a0abc000d, 48'hc191a87f035, 48'ha950795000c, 48'ha711b41ff74, 48'h9401b050001, 48'h83a0a770010, 48'h7043e1fffd5, 48'h7033e50ffcf, 48'h63c13cd0037, 48'h3dc31a9fff3, 48'h3db20561153, 48'h2a838c2ffec, 48'h15c0e940021, 48'h15b04010a93, 48'h3};
    //EXPECTED OUTPUT
    logic[`PWL_BRAM_DEPTH-1:0][`BATCH_SAMPLES-1:0][`SAMPLE_WIDTH-1:0] expected_batches;
    assign expected_batches = {0,{16'h097f, 16'h097f, 16'h097f, 16'h097f, 16'h097f, 16'h097f, 16'h097f, 16'h097f, 16'h097f, 16'h097f, 16'h097f, 16'h097f, 16'h0a20, 16'h0a3f, 16'h0a5e, 16'h0a7d, 16'h0a9c, 16'h0abb, 16'h0ada, 16'h0af9, 16'h0b18, 16'h0b37, 16'h0b56, 16'h0b75, 16'h0b94, 16'h0bb3, 16'h0bd2, 16'h0bf1, 16'h0c10, 16'h0c2f, 16'h0c4e, 16'h0c6d, 16'h0c8c, 16'h0cab, 16'h0cca, 16'h0ce9, 16'h0d08, 16'h0d27, 16'h0d46, 16'h0d65, 16'h0d84, 16'h0da3, 16'h0dc2, 16'h0de1, 16'h0e00, 16'h0e1f, 16'h0e3e, 16'h0e5d, 16'h0e7c, 16'h0e9b, 16'h0eba, 16'h0ed9, 16'h0ef8, 16'h0f17, 16'h0f36, 16'h0f55, 16'h0f74, 16'h0f93, 16'h0fb2, 16'h0fd1, 16'h0ff0, 16'h100f, 16'h102e, 16'h104d},
                                 {16'h106c, 16'h108b, 16'h10aa, 16'h10c9, 16'h10e8, 16'h1107, 16'h1126, 16'h1145, 16'h1164, 16'h1183, 16'h11a2, 16'h11c1, 16'h11e0, 16'h11ff, 16'h121e, 16'h123d, 16'h125c, 16'h127b, 16'h129a, 16'h12b9, 16'h12d8, 16'h12f7, 16'h1316, 16'h1335, 16'h1354, 16'h1373, 16'h1392, 16'h13b1, 16'h13d0, 16'h13ef, 16'h140e, 16'h142d, 16'h144c, 16'h146b, 16'h148a, 16'h14a9, 16'h14c8, 16'h14e7, 16'h1506, 16'h1525, 16'h1544, 16'h1563, 16'h1582, 16'h15a1, 16'h15c0, 16'h15df, 16'h15fe, 16'h161d, 16'h163c, 16'h165b, 16'h167a, 16'h1699, 16'h16b8, 16'h16d7, 16'h16f6, 16'h1715, 16'h1734, 16'h1753, 16'h1772, 16'h1791, 16'h17b0, 16'h17cf, 16'h17ee, 16'h180d},
                                 {16'h182c, 16'h184b, 16'h186a, 16'h1889, 16'h18a8, 16'h18c7, 16'h18e6, 16'h1905, 16'h1924, 16'h1943, 16'h1962, 16'h1981, 16'h19a0, 16'h19bf, 16'h19de, 16'h19fd, 16'h1a1c, 16'h1a3b, 16'h1a5a, 16'h1a79, 16'h1a98, 16'h1ab7, 16'h1ad6, 16'h1af5, 16'h1b14, 16'h1b33, 16'h1b52, 16'h1b71, 16'h1b90, 16'h1baf, 16'h1bce, 16'h1bed, 16'h1c0c, 16'h1c2b, 16'h1c4a, 16'h1c69, 16'h1c88, 16'h1ca7, 16'h1cc6, 16'h1ce5, 16'h1d04, 16'h1d23, 16'h1d42, 16'h1d61, 16'h1d80, 16'h1d9f, 16'h1dbe, 16'h1ddd, 16'h1dfc, 16'h1e1b, 16'h1e3a, 16'h1e59, 16'h1e78, 16'h1e97, 16'h1eb6, 16'h1ed5, 16'h1ef4, 16'h1f13, 16'h1f32, 16'h1f51, 16'h1f70, 16'h1f8f, 16'h1fae, 16'h1fcd},
                                 {16'h1fec, 16'h200b, 16'h202a, 16'h2049, 16'h2068, 16'h2087, 16'h20a6, 16'h20c5, 16'h20e4, 16'h2103, 16'h2122, 16'h2141, 16'h2160, 16'h217f, 16'h219e, 16'h21bd, 16'h21dc, 16'h21fb, 16'h221a, 16'h2239, 16'h2258, 16'h2277, 16'h2296, 16'h22b5, 16'h22d4, 16'h22f3, 16'h2312, 16'h2331, 16'h2350, 16'h236f, 16'h238e, 16'h23ad, 16'h23cc, 16'h23eb, 16'h240a, 16'h2429, 16'h2448, 16'h2467, 16'h2486, 16'h24a5, 16'h24c4, 16'h24e3, 16'h2502, 16'h2521, 16'h2540, 16'h255f, 16'h257e, 16'h259d, 16'h25bc, 16'h25db, 16'h25fa, 16'h2619, 16'h2638, 16'h2657, 16'h2676, 16'h2695, 16'h26b4, 16'h26d3, 16'h26f2, 16'h2711, 16'h2730, 16'h274f, 16'h276e, 16'h278d},
                                 {16'h27ac, 16'h27cb, 16'h27ea, 16'h2809, 16'h2828, 16'h2847, 16'h2866, 16'h2885, 16'h28a4, 16'h28c3, 16'h28e2, 16'h2901, 16'h2920, 16'h293f, 16'h295e, 16'h297d, 16'h299c, 16'h29bb, 16'h29da, 16'h29f9, 16'h2a18, 16'h2a37, 16'h2a56, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75},
                                 {16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75},
                                 {16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75},
                                 {16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75},
                                 {16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a75, 16'h2a76, 16'h2a77, 16'h2a78, 16'h2a79, 16'h2a7a, 16'h2a7b, 16'h2a7c, 16'h2a7d, 16'h2a7e, 16'h2a7f, 16'h2a80, 16'h2a81, 16'h2a82, 16'h2a83, 16'h2a84, 16'h2a85, 16'h2a86, 16'h2a87, 16'h2a88, 16'h2a89, 16'h2a8a, 16'h2a8b, 16'h2a8c, 16'h2a8d, 16'h2a78, 16'h2a54, 16'h2a30, 16'h2a0c, 16'h29e8, 16'h29c4, 16'h29a0, 16'h297c, 16'h2958, 16'h2934, 16'h2910, 16'h28ec, 16'h28c8, 16'h28a4, 16'h2880, 16'h285c, 16'h2838, 16'h2814, 16'h27f0, 16'h27cc, 16'h27a8, 16'h2784, 16'h2760, 16'h273c},
                                 {16'h2718, 16'h26f4, 16'h26d0, 16'h26ac, 16'h2688, 16'h2664, 16'h2640, 16'h261c, 16'h25f8, 16'h25d4, 16'h25b0, 16'h258c, 16'h2568, 16'h2544, 16'h2520, 16'h24fc, 16'h24d8, 16'h24b4, 16'h2490, 16'h246c, 16'h2448, 16'h2424, 16'h2400, 16'h23dc, 16'h23b8, 16'h2394, 16'h2370, 16'h234c, 16'h2328, 16'h2304, 16'h22e0, 16'h22bc, 16'h2298, 16'h2274, 16'h2250, 16'h222c, 16'h2208, 16'h21e4, 16'h21c0, 16'h219c, 16'h2178, 16'h2154, 16'h2130, 16'h210c, 16'h20e8, 16'h20c4, 16'h20a0, 16'h207c, 16'h2058, 16'h2034, 16'h2010, 16'h1fec, 16'h1fc8, 16'h1fa4, 16'h1f80, 16'h1f5c, 16'h1f38, 16'h1f14, 16'h1ef0, 16'h1ecc, 16'h1ea8, 16'h1e84, 16'h1e60, 16'h1e3c},
                                 {16'h1e18, 16'h1df4, 16'h1dd0, 16'h1dac, 16'h1d88, 16'h1d64, 16'h1d40, 16'h1d1c, 16'h1cf8, 16'h1cd4, 16'h1cb0, 16'h1c8c, 16'h1c68, 16'h1c44, 16'h1c20, 16'h1bfc, 16'h1bd8, 16'h1bb4, 16'h1b90, 16'h1b6c, 16'h1b48, 16'h1b24, 16'h1b00, 16'h1adc, 16'h1ab8, 16'h1a94, 16'h1a70, 16'h1a4c, 16'h1a28, 16'h1a04, 16'h19e0, 16'h19bc, 16'h1998, 16'h1974, 16'h1950, 16'h192c, 16'h1908, 16'h18e4, 16'h18c0, 16'h189c, 16'h1878, 16'h1854, 16'h1830, 16'h180c, 16'h17e8, 16'h17c4, 16'h17a0, 16'h177c, 16'h1758, 16'h1734, 16'h1710, 16'h16ec, 16'h16c8, 16'h16a4, 16'h1680, 16'h165c, 16'h1638, 16'h1614, 16'h15f0, 16'h15cc, 16'h15a8, 16'h1584, 16'h1560, 16'h153c},
                                 {16'h1518, 16'h14f4, 16'h14d0, 16'h14ac, 16'h1488, 16'h1464, 16'h1440, 16'h141c, 16'h13f8, 16'h13d4, 16'h13b0, 16'h138c, 16'h1368, 16'h1344, 16'h1320, 16'h12fc, 16'h12d8, 16'h12b4, 16'h1290, 16'h126c, 16'h1248, 16'h1224, 16'h1200, 16'h11dc, 16'h11b8, 16'h1194, 16'h1170, 16'h114c, 16'h1128, 16'h1104, 16'h10e0, 16'h10bc, 16'h1098, 16'h1074, 16'h1050, 16'h102c, 16'h1008, 16'h0fe4, 16'h0fc0, 16'h0f9c, 16'h0f78, 16'h0f54, 16'h0f30, 16'h0f0c, 16'h0ee8, 16'h0ec4, 16'h0ea0, 16'h0e7c, 16'h0e58, 16'h0e34, 16'h0e10, 16'h0dec, 16'h0dc8, 16'h0da4, 16'h0d80, 16'h0d5c, 16'h0d38, 16'h0d14, 16'h0cf0, 16'h0ccc, 16'h0ca8, 16'h0c84, 16'h0c60, 16'h0c3c},
                                 {16'h0c18, 16'h0bf4, 16'h0bd0, 16'h0bac, 16'h0b88, 16'h0b64, 16'h0b40, 16'h0b1c, 16'h0af8, 16'h0ad4, 16'h0ab0, 16'h0a8c, 16'h0a68, 16'h0a44, 16'h0a20, 16'h09fc, 16'h09d8, 16'h09b4, 16'h0990, 16'h096c, 16'h0948, 16'h0924, 16'h0900, 16'h08dc, 16'h08b8, 16'h0894, 16'h0870, 16'h084c, 16'h0828, 16'h0804, 16'h07e0, 16'h07bc, 16'h0798, 16'h0774, 16'h0750, 16'h072c, 16'h0708, 16'h06e4, 16'h06c0, 16'h069c, 16'h0678, 16'h0654, 16'h0630, 16'h060c, 16'h05e8, 16'h05c4, 16'h05a0, 16'h057c, 16'h0558, 16'h0534, 16'h0510, 16'h04ec, 16'h04c8, 16'h04a4, 16'h0480, 16'h045c, 16'h0438, 16'h0414, 16'h0414, 16'h0414, 16'h0414, 16'h0414, 16'h0414, 16'h0414},
                                 {16'h0414, 16'h0414, 16'h0414, 16'h0414, 16'h0414, 16'h0414, 16'h0413, 16'h0412, 16'h0411, 16'h0410, 16'h040f, 16'h040e, 16'h040d, 16'h040c, 16'h040b, 16'h040a, 16'h0409, 16'h0408, 16'h0407, 16'h0406, 16'h0405, 16'h0404, 16'h0403, 16'h0402, 16'h0401, 16'h0400, 16'h03ff, 16'h03fe, 16'h03fd, 16'h03fc, 16'h03fb, 16'h03fa, 16'h03f9, 16'h03f8, 16'h03f7, 16'h03f6, 16'h03f5, 16'h03f4, 16'h03f3, 16'h03f2, 16'h03f1, 16'h03f0, 16'h03ef, 16'h03ee, 16'h03ed, 16'h03ec, 16'h03eb, 16'h03ea, 16'h03e9, 16'h03e8, 16'h03e7, 16'h03e6, 16'h03e5, 16'h03e4, 16'h03e3, 16'h03e2, 16'h03e1, 16'h03e0, 16'h03df, 16'h03de, 16'h03dd, 16'h03dc, 16'h03db, 16'h03da},
                                 {16'h03d9, 16'h03d8, 16'h03d7, 16'h03d6, 16'h03d5, 16'h03d4, 16'h03d3, 16'h03d2, 16'h03d1, 16'h03d0, 16'h03cf, 16'h03ce, 16'h03cd, 16'h03cc, 16'h03cb, 16'h03ca, 16'h03c9, 16'h03c8, 16'h03c7, 16'h03c6, 16'h03c5, 16'h03c4, 16'h03c3, 16'h03c2, 16'h03c1, 16'h03c0, 16'h03bf, 16'h03be, 16'h03bd, 16'h03bc, 16'h03bb, 16'h03ba, 16'h03b9, 16'h03b8, 16'h03b7, 16'h03b6, 16'h03b5, 16'h03b4, 16'h03b3, 16'h03b2, 16'h03b1, 16'h03b0, 16'h03af, 16'h03ae, 16'h03ad, 16'h03ac, 16'h03ab, 16'h03aa, 16'h03a9, 16'h03a8, 16'h03a7, 16'h03a6, 16'h03a5, 16'h03a4, 16'h03a3, 16'h03a2, 16'h03a1, 16'h03a0, 16'h039f, 16'h039e, 16'h039d, 16'h039c, 16'h039b, 16'h039a},
                                 {16'h0399, 16'h0398, 16'h0397, 16'h0396, 16'h0395, 16'h0394, 16'h0393, 16'h0392, 16'h0391, 16'h0390, 16'h038f, 16'h038e, 16'h038d, 16'h038c, 16'h038b, 16'h038a, 16'h0389, 16'h0388, 16'h0387, 16'h0386, 16'h0385, 16'h0384, 16'h0383, 16'h0382, 16'h0381, 16'h0380, 16'h037f, 16'h037e, 16'h037d, 16'h037c, 16'h037b, 16'h037a, 16'h0379, 16'h0378, 16'h0377, 16'h0376, 16'h0375, 16'h0374, 16'h0373, 16'h0372, 16'h0371, 16'h0370, 16'h036f, 16'h036e, 16'h036d, 16'h036c, 16'h036b, 16'h036a, 16'h0369, 16'h0368, 16'h0367, 16'h0366, 16'h0365, 16'h0364, 16'h0363, 16'h0362, 16'h0361, 16'h0360, 16'h035f, 16'h035e, 16'h035d, 16'h035c, 16'h035b, 16'h035a},
                                 {16'h0359, 16'h0358, 16'h0357, 16'h0356, 16'h0355, 16'h0354, 16'h0353, 16'h0352, 16'h0351, 16'h0350, 16'h034f, 16'h034e, 16'h034d, 16'h034c, 16'h034b, 16'h034a, 16'h0349, 16'h0348, 16'h0347, 16'h0346, 16'h0345, 16'h0344, 16'h0343, 16'h0342, 16'h0341, 16'h0340, 16'h033f, 16'h033e, 16'h033d, 16'h033c, 16'h033b, 16'h033a, 16'h0339, 16'h0338, 16'h0337, 16'h0336, 16'h0335, 16'h0334, 16'h0333, 16'h0332, 16'h0331, 16'h0330, 16'h032f, 16'h032e, 16'h032d, 16'h032c, 16'h032b, 16'h032a, 16'h0329, 16'h0328, 16'h0327, 16'h0326, 16'h0325, 16'h0324, 16'h0323, 16'h0322, 16'h0321, 16'h0320, 16'h031f, 16'h031e, 16'h031d, 16'h031c, 16'h031b, 16'h031a},
                                 {16'h0319, 16'h0318, 16'h0317, 16'h0316, 16'h0315, 16'h0314, 16'h0313, 16'h0312, 16'h0311, 16'h0310, 16'h030f, 16'h030e, 16'h030d, 16'h030c, 16'h030b, 16'h030a, 16'h0309, 16'h0308, 16'h0307, 16'h0306, 16'h0305, 16'h0304, 16'h0303, 16'h0302, 16'h0301, 16'h0300, 16'h02ff, 16'h02fe, 16'h02fd, 16'h02fc, 16'h02fb, 16'h02fa, 16'h02f9, 16'h02f8, 16'h02f7, 16'h02f6, 16'h02f5, 16'h02f4, 16'h02f3, 16'h02f2, 16'h02f1, 16'h02f0, 16'h02ef, 16'h02ee, 16'h02ed, 16'h02ec, 16'h02eb, 16'h02ea, 16'h02e9, 16'h02e8, 16'h02e7, 16'h02e6, 16'h02e5, 16'h02e4, 16'h02e3, 16'h02e2, 16'h02e1, 16'h02e0, 16'h02df, 16'h02de, 16'h02dd, 16'h02dc, 16'h02db, 16'h02da},
                                 {16'h02d9, 16'h02d8, 16'h02d7, 16'h02d6, 16'h02d5, 16'h02d4, 16'h02d3, 16'h02d2, 16'h02d1, 16'h02d0, 16'h02cf, 16'h02ce, 16'h02cd, 16'h02cc, 16'h02cb, 16'h02ca, 16'h02c9, 16'h02c8, 16'h02c7, 16'h02c6, 16'h02c5, 16'h02c4, 16'h02c3, 16'h02c2, 16'h02c1, 16'h02c0, 16'h02bf, 16'h02be, 16'h02bd, 16'h02bc, 16'h02bb, 16'h02ba, 16'h02b9, 16'h02b8, 16'h02b7, 16'h02b6, 16'h02b5, 16'h02b4, 16'h02b3, 16'h02b2, 16'h02b1, 16'h02b0, 16'h02af, 16'h02ae, 16'h02ad, 16'h02ac, 16'h02ab, 16'h02aa, 16'h02a9, 16'h02a8, 16'h02a7, 16'h02a6, 16'h02a5, 16'h02a4, 16'h02a3, 16'h02a2, 16'h02a1, 16'h02a0, 16'h029f, 16'h029e, 16'h029d, 16'h029c, 16'h029b, 16'h029a},
                                 {16'h0299, 16'h0298, 16'h0297, 16'h0296, 16'h0295, 16'h0294, 16'h0293, 16'h0292, 16'h0291, 16'h0290, 16'h028f, 16'h028e, 16'h028d, 16'h028c, 16'h028b, 16'h028a, 16'h0289, 16'h0288, 16'h0287, 16'h0286, 16'h0285, 16'h0284, 16'h0283, 16'h0282, 16'h0281, 16'h0280, 16'h027f, 16'h027e, 16'h027d, 16'h027c, 16'h027b, 16'h027a, 16'h0279, 16'h0278, 16'h0277, 16'h0276, 16'h0275, 16'h0274, 16'h0273, 16'h0272, 16'h0271, 16'h0270, 16'h02b8, 16'h031f, 16'h0386, 16'h03ed, 16'h0454, 16'h04bb, 16'h0522, 16'h0589, 16'h05f0, 16'h0657, 16'h06be, 16'h0725, 16'h078c, 16'h07f3, 16'h085a, 16'h08c1, 16'h0928, 16'h098f, 16'h09f6, 16'h0a5d, 16'h0ac4, 16'h0b2b},
                                 {16'h0b92, 16'h0bf9, 16'h0c60, 16'h0cc7, 16'h0d2e, 16'h0d95, 16'h0dfc, 16'h0e63, 16'h0eca, 16'h0f31, 16'h0f98, 16'h0fff, 16'h1066, 16'h10cd, 16'h1134, 16'h119b, 16'h1202, 16'h1269, 16'h12d0, 16'h1337, 16'h139e, 16'h1405, 16'h146c, 16'h14d3, 16'h153a, 16'h15a1, 16'h1608, 16'h166f, 16'h16d6, 16'h173d, 16'h17a4, 16'h180b, 16'h1872, 16'h18d9, 16'h1940, 16'h19a7, 16'h1a0e, 16'h1a75, 16'h1adc, 16'h1b43, 16'h1baa, 16'h1c11, 16'h1c78, 16'h1cdf, 16'h1d46, 16'h1dad, 16'h1e14, 16'h1e7b, 16'h1ee2, 16'h1f49, 16'h1fb0, 16'h2017, 16'h207e, 16'h20e5, 16'h214c, 16'h21b3, 16'h221a, 16'h2281, 16'h22e8, 16'h234f, 16'h23b6, 16'h241d, 16'h2484, 16'h24eb},
                                 {16'h2552, 16'h25b9, 16'h2620, 16'h2687, 16'h26ee, 16'h2755, 16'h27bc, 16'h2823, 16'h288a, 16'h28f1, 16'h2958, 16'h29bf, 16'h2a26, 16'h2a8d, 16'h2af4, 16'h2b5b, 16'h2bc2, 16'h2c29, 16'h2c90, 16'h2cf7, 16'h2d5e, 16'h2dc5, 16'h2e2c, 16'h2e93, 16'h2efa, 16'h2f61, 16'h2fc8, 16'h302f, 16'h3096, 16'h30fd, 16'h3164, 16'h31cb, 16'h3232, 16'h3299, 16'h3300, 16'h3367, 16'h33ce, 16'h3435, 16'h349c, 16'h3503, 16'h356a, 16'h35d1, 16'h3638, 16'h369f, 16'h3706, 16'h376d, 16'h37d4, 16'h383b, 16'h38a2, 16'h3909, 16'h3970, 16'h39d7, 16'h3a3e, 16'h3a4f, 16'h3a58, 16'h3a61, 16'h3a6a, 16'h3a73, 16'h3a7c, 16'h3a85, 16'h3a8e, 16'h3a97, 16'h3aa0, 16'h3aa9},
                                 {16'h3ab2, 16'h3abb, 16'h3ac4, 16'h3acd, 16'h3ad6, 16'h3adf, 16'h3ae8, 16'h3af1, 16'h3afa, 16'h3b03, 16'h3b0c, 16'h3b15, 16'h3b1e, 16'h3b27, 16'h3b30, 16'h3b39, 16'h3b42, 16'h3b4b, 16'h3b54, 16'h3b5d, 16'h3b66, 16'h3b6f, 16'h3b78, 16'h3b81, 16'h3b8a, 16'h3b93, 16'h3b9c, 16'h3ba5, 16'h3bae, 16'h3bb7, 16'h3bc0, 16'h3bc9, 16'h3bd2, 16'h3bdb, 16'h3be4, 16'h3bed, 16'h3bf6, 16'h3bff, 16'h3c08, 16'h3c11, 16'h3c1a, 16'h3c23, 16'h3c2c, 16'h3c35, 16'h3c3e, 16'h3c47, 16'h3c50, 16'h3c59, 16'h3c62, 16'h3c6b, 16'h3c74, 16'h3c7d, 16'h3c86, 16'h3c8f, 16'h3c98, 16'h3ca1, 16'h3caa, 16'h3cb3, 16'h3cbc, 16'h3cc5, 16'h3cce, 16'h3cd7, 16'h3ce0, 16'h3ce9},
                                 {16'h3cf2, 16'h3cfb, 16'h3d04, 16'h3d0d, 16'h3d16, 16'h3d1f, 16'h3d28, 16'h3d31, 16'h3d3a, 16'h3d43, 16'h3d4c, 16'h3d55, 16'h3d5e, 16'h3d67, 16'h3d70, 16'h3d79, 16'h3d53, 16'h3d3d, 16'h3d27, 16'h3d11, 16'h3cfb, 16'h3ce5, 16'h3ccf, 16'h3cb9, 16'h3ca3, 16'h3c8d, 16'h3c77, 16'h3c61, 16'h3c4b, 16'h3c35, 16'h3c1f, 16'h3c09, 16'h3bf3, 16'h3bdd, 16'h3bc7, 16'h3bb1, 16'h3b9b, 16'h3b85, 16'h3b6f, 16'h3b59, 16'h3b43, 16'h3b2d, 16'h3b17, 16'h3b01, 16'h3aeb, 16'h3ad5, 16'h3abf, 16'h3aa9, 16'h3a93, 16'h3a7d, 16'h3a67, 16'h3a51, 16'h3a3b, 16'h3a25, 16'h3a0f, 16'h39f9, 16'h39e3, 16'h39cd, 16'h39b7, 16'h39a1, 16'h398b, 16'h3975, 16'h395f, 16'h3949},
                                 {16'h3933, 16'h391d, 16'h3907, 16'h38f1, 16'h38db, 16'h38c5, 16'h38af, 16'h3899, 16'h3883, 16'h386d, 16'h3857, 16'h3841, 16'h382b, 16'h3815, 16'h37ff, 16'h37e9, 16'h37d3, 16'h37bd, 16'h37a7, 16'h3791, 16'h377b, 16'h3765, 16'h374f, 16'h3739, 16'h3723, 16'h370d, 16'h36f7, 16'h36e1, 16'h36cb, 16'h36b5, 16'h369f, 16'h3689, 16'h3673, 16'h365d, 16'h3647, 16'h3631, 16'h361b, 16'h3605, 16'h35ef, 16'h35d9, 16'h35c3, 16'h35ad, 16'h3597, 16'h3581, 16'h356b, 16'h3555, 16'h353f, 16'h3529, 16'h3513, 16'h34fd, 16'h34e7, 16'h34d1, 16'h34bb, 16'h34a5, 16'h348f, 16'h3479, 16'h3463, 16'h344d, 16'h3437, 16'h3421, 16'h340b, 16'h33f5, 16'h33df, 16'h33c9},
                                 {16'h33b3, 16'h339d, 16'h3387, 16'h3371, 16'h335b, 16'h3345, 16'h332f, 16'h3319, 16'h3303, 16'h32ed, 16'h32d7, 16'h32c1, 16'h32ab, 16'h3295, 16'h327f, 16'h3269, 16'h3253, 16'h323d, 16'h3227, 16'h3211, 16'h31fb, 16'h31e5, 16'h31cf, 16'h31b9, 16'h31a3, 16'h318d, 16'h3177, 16'h3161, 16'h314b, 16'h3135, 16'h311f, 16'h3109, 16'h30f3, 16'h30dd, 16'h30c7, 16'h30b1, 16'h309b, 16'h3085, 16'h306f, 16'h3059, 16'h3043, 16'h302d, 16'h3017, 16'h3001, 16'h2feb, 16'h2fd5, 16'h2fbf, 16'h2fa9, 16'h2f93, 16'h2f7d, 16'h2f67, 16'h2f51, 16'h2f3b, 16'h2f25, 16'h2f0f, 16'h2ef9, 16'h2ee3, 16'h2ecd, 16'h2eb7, 16'h2ea1, 16'h2e8b, 16'h2e75, 16'h2e5f, 16'h2e49},
                                 {16'h2e33, 16'h2e1d, 16'h2e07, 16'h2df1, 16'h2ddb, 16'h2dc5, 16'h2daf, 16'h2d99, 16'h2d83, 16'h2d6d, 16'h2d57, 16'h2d41, 16'h2d2b, 16'h2d15, 16'h2cff, 16'h2ce9, 16'h2cd3, 16'h2cbd, 16'h2ca7, 16'h2c91, 16'h2c7b, 16'h2c65, 16'h2c4f, 16'h2c39, 16'h2c23, 16'h2c0d, 16'h2bf7, 16'h2be1, 16'h2bcb, 16'h2bb5, 16'h2b9f, 16'h2b89, 16'h2b73, 16'h2b5d, 16'h2b47, 16'h2b31, 16'h2b1b, 16'h2b05, 16'h2aef, 16'h2ad9, 16'h2ac3, 16'h2aad, 16'h2a97, 16'h2a81, 16'h2a6b, 16'h2a55, 16'h2a3f, 16'h2a29, 16'h2a13, 16'h29fd, 16'h29e7, 16'h29d1, 16'h29bb, 16'h29a5, 16'h298f, 16'h2979, 16'h2963, 16'h294d, 16'h2937, 16'h2921, 16'h290b, 16'h28f5, 16'h28df, 16'h28c9},
                                 {16'h28b3, 16'h289d, 16'h2887, 16'h2871, 16'h285b, 16'h2845, 16'h282f, 16'h2819, 16'h2803, 16'h27ed, 16'h27d7, 16'h27c1, 16'h27ab, 16'h2795, 16'h277f, 16'h2769, 16'h2753, 16'h273d, 16'h2727, 16'h2711, 16'h26fb, 16'h26e5, 16'h26cf, 16'h26b9, 16'h26a3, 16'h268d, 16'h2677, 16'h2661, 16'h264b, 16'h2635, 16'h261f, 16'h2609, 16'h25f3, 16'h25dd, 16'h25c7, 16'h25b1, 16'h259b, 16'h2585, 16'h256f, 16'h2559, 16'h2543, 16'h252d, 16'h2517, 16'h2501, 16'h24eb, 16'h24d5, 16'h24bf, 16'h24a9, 16'h2493, 16'h247d, 16'h2467, 16'h2451, 16'h243b, 16'h2425, 16'h240f, 16'h23f9, 16'h23e3, 16'h23cd, 16'h23b7, 16'h23a1, 16'h238b, 16'h2375, 16'h235f, 16'h2349},
                                 {16'h2333, 16'h231d, 16'h2307, 16'h22f1, 16'h22db, 16'h22c5, 16'h22af, 16'h2299, 16'h2283, 16'h226d, 16'h2257, 16'h2241, 16'h222b, 16'h2215, 16'h21ff, 16'h21e9, 16'h21d3, 16'h21bd, 16'h21a7, 16'h2191, 16'h217b, 16'h2165, 16'h214f, 16'h2139, 16'h2123, 16'h210d, 16'h20f7, 16'h20e1, 16'h20cb, 16'h20b5, 16'h209f, 16'h2089, 16'h2073, 16'h205d, 16'h2047, 16'h2031, 16'h201b, 16'h2005, 16'h1fef, 16'h1fd9, 16'h1fc3, 16'h1fad, 16'h1f97, 16'h1f81, 16'h1f6b, 16'h1f55, 16'h1f3f, 16'h1f29, 16'h1f13, 16'h1efd, 16'h1ee7, 16'h1ed1, 16'h1ebb, 16'h1ea5, 16'h1e8f, 16'h1e79, 16'h1e63, 16'h1e4d, 16'h1e37, 16'h1e21, 16'h1e0b, 16'h1df5, 16'h1ddf, 16'h1dc9},
                                 {16'h1db3, 16'h1d9d, 16'h1d87, 16'h1d71, 16'h1d5b, 16'h1d45, 16'h1d2f, 16'h1d19, 16'h1d03, 16'h1d57, 16'h1d78, 16'h1d99, 16'h1dba, 16'h1ddb, 16'h1dfc, 16'h1e1d, 16'h1e3e, 16'h1e5f, 16'h1e80, 16'h1ea1, 16'h1ec2, 16'h1ee3, 16'h1f04, 16'h1f25, 16'h1f46, 16'h1f67, 16'h1f88, 16'h1fa9, 16'h1fca, 16'h1feb, 16'h200c, 16'h202d, 16'h204e, 16'h206f, 16'h2090, 16'h20b1, 16'h20d2, 16'h20f3, 16'h2114, 16'h2135, 16'h2156, 16'h2177, 16'h2198, 16'h21b9, 16'h21da, 16'h21fb, 16'h221c, 16'h223d, 16'h225e, 16'h227f, 16'h22a0, 16'h22c1, 16'h22e2, 16'h2303, 16'h2324, 16'h2345, 16'h2366, 16'h2387, 16'h23a8, 16'h23c9, 16'h23ea, 16'h240b, 16'h242c, 16'h244d},
                                 {16'h246e, 16'h248f, 16'h24b0, 16'h24d1, 16'h24f2, 16'h2513, 16'h2534, 16'h2555, 16'h2576, 16'h2597, 16'h25b8, 16'h25d9, 16'h25fa, 16'h261b, 16'h263c, 16'h265d, 16'h267e, 16'h269f, 16'h26c0, 16'h26e1, 16'h2702, 16'h2723, 16'h2744, 16'h2765, 16'h2786, 16'h27a7, 16'h27c8, 16'h27e9, 16'h280a, 16'h282b, 16'h284c, 16'h286d, 16'h288e, 16'h28af, 16'h28d0, 16'h28f1, 16'h2912, 16'h2933, 16'h2954, 16'h2975, 16'h2996, 16'h29b7, 16'h29d8, 16'h29f9, 16'h2a1a, 16'h2a3b, 16'h2a5c, 16'h2a7d, 16'h2a9e, 16'h2abf, 16'h2ae0, 16'h2b01, 16'h2b22, 16'h2b43, 16'h2b64, 16'h2b85, 16'h2ba6, 16'h2bc7, 16'h2be8, 16'h2c09, 16'h2c2a, 16'h2c4b, 16'h2c6c, 16'h2c8d},
                                 {16'h2cae, 16'h2ccf, 16'h2cf0, 16'h2d11, 16'h2d32, 16'h2d53, 16'h2d74, 16'h2d95, 16'h2db6, 16'h2dd7, 16'h2df8, 16'h2e19, 16'h2e3a, 16'h2e5b, 16'h2e7c, 16'h2e9d, 16'h2ebe, 16'h2edf, 16'h2f00, 16'h2f21, 16'h2f42, 16'h2f63, 16'h2f84, 16'h2fa5, 16'h2fc6, 16'h2fe7, 16'h3008, 16'h3029, 16'h304a, 16'h306b, 16'h308c, 16'h30ad, 16'h30ce, 16'h30ef, 16'h3110, 16'h3131, 16'h3152, 16'h3173, 16'h3194, 16'h31b5, 16'h31d6, 16'h31f7, 16'h3218, 16'h3239, 16'h325a, 16'h327b, 16'h329c, 16'h32bd, 16'h32de, 16'h32ff, 16'h3320, 16'h3341, 16'h3362, 16'h3383, 16'h33a4, 16'h33c5, 16'h33e6, 16'h3407, 16'h3428, 16'h3449, 16'h346a, 16'h342d, 16'h3413, 16'h33f9},
                                 {16'h33df, 16'h33c5, 16'h33ab, 16'h3391, 16'h3377, 16'h335d, 16'h3343, 16'h3329, 16'h330f, 16'h32f5, 16'h32db, 16'h32c1, 16'h32a7, 16'h328d, 16'h3273, 16'h3259, 16'h323f, 16'h3225, 16'h320b, 16'h31f1, 16'h31d7, 16'h31bd, 16'h31a3, 16'h3189, 16'h316f, 16'h3155, 16'h313b, 16'h3121, 16'h3107, 16'h30ed, 16'h30d3, 16'h30b9, 16'h309f, 16'h3085, 16'h306b, 16'h3051, 16'h3037, 16'h301d, 16'h3003, 16'h2fe9, 16'h2fcf, 16'h2fb5, 16'h2f9b, 16'h2f81, 16'h2f67, 16'h2f4d, 16'h2f33, 16'h2f19, 16'h2eff, 16'h2ee5, 16'h2ecb, 16'h2eb1, 16'h2e97, 16'h2e7d, 16'h2e63, 16'h2e49, 16'h2e2f, 16'h2e15, 16'h2dfb, 16'h2de1, 16'h2dc7, 16'h2dad, 16'h2d93, 16'h2d79},
                                 {16'h2d5f, 16'h2d45, 16'h2d2b, 16'h2d11, 16'h2cf7, 16'h2cdd, 16'h2cc3, 16'h2ca9, 16'h2c8f, 16'h2c75, 16'h2c5b, 16'h2c41, 16'h2c27, 16'h2c0d, 16'h2bf3, 16'h2bd9, 16'h2bbf, 16'h2ba5, 16'h2b8b, 16'h2b71, 16'h2b57, 16'h2b3d, 16'h2b23, 16'h2b09, 16'h2aef, 16'h2ad5, 16'h2abb, 16'h2aa1, 16'h2a87, 16'h2a6d, 16'h2a53, 16'h2a39, 16'h2a1f, 16'h2a05, 16'h29eb, 16'h29d1, 16'h29b7, 16'h299d, 16'h2983, 16'h2969, 16'h294f, 16'h2935, 16'h291b, 16'h2901, 16'h28e7, 16'h28cd, 16'h28b3, 16'h2899, 16'h287f, 16'h2865, 16'h284b, 16'h2831, 16'h2817, 16'h27fd, 16'h27e3, 16'h27c9, 16'h27af, 16'h2795, 16'h277b, 16'h2761, 16'h2747, 16'h272d, 16'h2713, 16'h26f9},
                                 {16'h26df, 16'h26c5, 16'h26ab, 16'h2691, 16'h2677, 16'h265d, 16'h2643, 16'h2629, 16'h260f, 16'h25f5, 16'h25db, 16'h25c1, 16'h25a7, 16'h258d, 16'h2573, 16'h2559, 16'h253f, 16'h2525, 16'h250b, 16'h24f1, 16'h24d7, 16'h24bd, 16'h24a3, 16'h2489, 16'h246f, 16'h2455, 16'h243b, 16'h2421, 16'h2407, 16'h23ed, 16'h23d3, 16'h23b9, 16'h239f, 16'h2385, 16'h236b, 16'h2351, 16'h2337, 16'h231d, 16'h2303, 16'h22e9, 16'h22cf, 16'h22b5, 16'h229b, 16'h2281, 16'h2267, 16'h224d, 16'h2233, 16'h2219, 16'h21ff, 16'h21e5, 16'h21cb, 16'h21b1, 16'h2197, 16'h217d, 16'h2163, 16'h2149, 16'h212f, 16'h2115, 16'h20fb, 16'h20e1, 16'h20c7, 16'h20ad, 16'h2093, 16'h2079},
                                 {16'h205f, 16'h2045, 16'h202b, 16'h2011, 16'h1ff7, 16'h1fdd, 16'h1fc3, 16'h1fa9, 16'h1f8f, 16'h1f75, 16'h1f5b, 16'h1f41, 16'h1f27, 16'h1f0d, 16'h1ef3, 16'h1ed9, 16'h1ebf, 16'h1ea5, 16'h1e8b, 16'h1e71, 16'h1e57, 16'h1e3d, 16'h1e23, 16'h1e09, 16'h1def, 16'h1dd5, 16'h1dbb, 16'h1da1, 16'h1d87, 16'h1d6d, 16'h1d53, 16'h1d39, 16'h1d1f, 16'h1d05, 16'h1ceb, 16'h1cd1, 16'h1cb7, 16'h1c9d, 16'h1c83, 16'h1c69, 16'h1c4f, 16'h1c35, 16'h1c1b, 16'h1c01, 16'h1be7, 16'h1bcd, 16'h1bb3, 16'h1b99, 16'h1b7f, 16'h1b65, 16'h1b4b, 16'h1b31, 16'h1b17, 16'h1afd, 16'h1ae3, 16'h1ac9, 16'h1aaf, 16'h1a95, 16'h1a7b, 16'h1a61, 16'h1a47, 16'h1a2d, 16'h1a13, 16'h19f9},
                                 {16'h19df, 16'h19c5, 16'h19ab, 16'h1991, 16'h1977, 16'h195d, 16'h1943, 16'h1929, 16'h190f, 16'h18f5, 16'h18db, 16'h18c1, 16'h18a7, 16'h188d, 16'h1873, 16'h1859, 16'h183f, 16'h1825, 16'h180b, 16'h17f1, 16'h17d7, 16'h17bd, 16'h17a3, 16'h1789, 16'h176f, 16'h1755, 16'h173b, 16'h1721, 16'h1707, 16'h16ed, 16'h16d3, 16'h16b9, 16'h169f, 16'h1685, 16'h166b, 16'h1651, 16'h1637, 16'h161d, 16'h1603, 16'h15e9, 16'h15cf, 16'h15b5, 16'h159b, 16'h1581, 16'h1567, 16'h154d, 16'h1533, 16'h1519, 16'h14ff, 16'h14e5, 16'h14cb, 16'h14b1, 16'h1497, 16'h147d, 16'h1463, 16'h1449, 16'h142f, 16'h1415, 16'h13fb, 16'h13e1, 16'h13c7, 16'h13ad, 16'h1393, 16'h1379},
                                 {16'h135f, 16'h1345, 16'h132b, 16'h1311, 16'h12f7, 16'h12dd, 16'h12c3, 16'h12a9, 16'h128f, 16'h1275, 16'h125b, 16'h1241, 16'h1227, 16'h120d, 16'h11f3, 16'h11d9, 16'h11bf, 16'h11a5, 16'h118b, 16'h1171, 16'h1157, 16'h113d, 16'h1123, 16'h1109, 16'h10ef, 16'h10d5, 16'h10bb, 16'h10a1, 16'h1087, 16'h106d, 16'h1053, 16'h1039, 16'h101f, 16'h1005, 16'h0feb, 16'h0fd1, 16'h0fb7, 16'h0f9d, 16'h0f83, 16'h0f69, 16'h0f4f, 16'h0f35, 16'h0f1b, 16'h0f01, 16'h0ee7, 16'h0ecd, 16'h0eb3, 16'h0e99, 16'h0e7f, 16'h0e65, 16'h0e4b, 16'h0e31, 16'h0e17, 16'h0dfd, 16'h0de3, 16'h0dc9, 16'h0daf, 16'h0d95, 16'h0d7b, 16'h0d61, 16'h0d47, 16'h0d2d, 16'h0d13, 16'h0cf9},
                                 {16'h0cdf, 16'h0cc5, 16'h0cab, 16'h0c91, 16'h0c77, 16'h0c5d, 16'h0c43, 16'h0c29, 16'h0c0f, 16'h0bf5, 16'h0bdb, 16'h0bc1, 16'h0ba7, 16'h0b8d, 16'h0b73, 16'h0b59, 16'h0b3f, 16'h0b25, 16'h0b0b, 16'h0af1, 16'h0ad7, 16'h0abd, 16'h0aa3, 16'h0a89, 16'h0a6f, 16'h0a55, 16'h0a3b, 16'h0a21, 16'h0a07, 16'h09ed, 16'h09d3, 16'h09b9, 16'h099f, 16'h0985, 16'h096b, 16'h0951, 16'h0937, 16'h091d, 16'h0903, 16'h08e9, 16'h08cf, 16'h08b5, 16'h089b, 16'h0881, 16'h0867, 16'h084d, 16'h0833, 16'h0819, 16'h07ff, 16'h07e5, 16'h07cb, 16'h07b1, 16'h0797, 16'h077d, 16'h0763, 16'h0749, 16'h072f, 16'h0715, 16'h06fb, 16'h06e1, 16'h06c7, 16'h06ad, 16'h0693, 16'h0679},
                                 {16'h065f, 16'h0645, 16'h062b, 16'h0611, 16'h05f7, 16'h05dd, 16'h05c3, 16'h05a9, 16'h058f, 16'h0575, 16'h055b, 16'h0541, 16'h0527, 16'h050d, 16'h04f3, 16'h04de, 16'h04d8, 16'h04d2, 16'h04cc, 16'h04c6, 16'h04c0, 16'h04ba, 16'h04b4, 16'h04ae, 16'h04a8, 16'h04a2, 16'h049c, 16'h0496, 16'h0490, 16'h048a, 16'h0484, 16'h047e, 16'h0478, 16'h0472, 16'h046c, 16'h0466, 16'h0460, 16'h045a, 16'h0454, 16'h044e, 16'h0448, 16'h0442, 16'h043c, 16'h0436, 16'h0430, 16'h042a, 16'h0424, 16'h041e, 16'h0418, 16'h0412, 16'h040c, 16'h042d, 16'h0440, 16'h0453, 16'h0466, 16'h0479, 16'h048c, 16'h049f, 16'h04b2, 16'h04c5, 16'h04d8, 16'h04eb, 16'h04fe, 16'h0511},
                                 {16'h0524, 16'h0537, 16'h054a, 16'h055d, 16'h0570, 16'h0583, 16'h0596, 16'h05a9, 16'h05bc, 16'h05cf, 16'h05e2, 16'h05f5, 16'h0608, 16'h061b, 16'h062e, 16'h0641, 16'h0654, 16'h0667, 16'h067a, 16'h068d, 16'h06a0, 16'h06b3, 16'h06c6, 16'h06d9, 16'h06ec, 16'h06ff, 16'h0712, 16'h0725, 16'h0738, 16'h074b, 16'h075e, 16'h0771, 16'h0784, 16'h0797, 16'h07aa, 16'h07bd, 16'h07d0, 16'h07e3, 16'h07f6, 16'h0809, 16'h081c, 16'h082f, 16'h0842, 16'h0855, 16'h0868, 16'h087b, 16'h088e, 16'h08a1, 16'h08b4, 16'h08c7, 16'h08da, 16'h08ed, 16'h0900, 16'h0913, 16'h0926, 16'h0939, 16'h094c, 16'h095f, 16'h0972, 16'h0985, 16'h0998, 16'h09ab, 16'h09be, 16'h09d1},
                                 {16'h09e4, 16'h09f7, 16'h0a0a, 16'h0a1d, 16'h0a30, 16'h0a43, 16'h0a56, 16'h0a69, 16'h0a7c, 16'h0a8f, 16'h0aa2, 16'h0ab5, 16'h0ac8, 16'h0adb, 16'h0aee, 16'h0b01, 16'h0b14, 16'h0b27, 16'h0b3a, 16'h0b4d, 16'h0b60, 16'h0b73, 16'h0b86, 16'h0b99, 16'h0bac, 16'h0bbf, 16'h0bd2, 16'h0be5, 16'h0bf8, 16'h0c0b, 16'h0c1e, 16'h0c31, 16'h0c44, 16'h0c57, 16'h0c6a, 16'h0c7d, 16'h0c90, 16'h0ca3, 16'h0cb6, 16'h0cc9, 16'h0cdc, 16'h0cef, 16'h0d02, 16'h0d15, 16'h0d28, 16'h0d3b, 16'h0d4e, 16'h0d61, 16'h0d74, 16'h0d87, 16'h0d9a, 16'h0dad, 16'h0dc0, 16'h0dd3, 16'h0de6, 16'h0df9, 16'h0e0c, 16'h0e1f, 16'h0e32, 16'h0e45, 16'h0e58, 16'h0e6b, 16'h0e7e, 16'h0e91},
                                 {16'h0ea4, 16'h0eb7, 16'h0eca, 16'h0edd, 16'h0ef0, 16'h0f03, 16'h0f16, 16'h0f29, 16'h0f3c, 16'h0f4f, 16'h0f62, 16'h0f75, 16'h0f88, 16'h0f9b, 16'h0fae, 16'h0fc1, 16'h0fd4, 16'h0fe7, 16'h0ffa, 16'h100d, 16'h1020, 16'h1033, 16'h1046, 16'h1059, 16'h106c, 16'h107f, 16'h1092, 16'h10a5, 16'h10b8, 16'h10cb, 16'h10de, 16'h10f1, 16'h1104, 16'h1117, 16'h112a, 16'h113d, 16'h1150, 16'h1163, 16'h1176, 16'h1189, 16'h119c, 16'h11af, 16'h11c2, 16'h11d5, 16'h11e8, 16'h11fb, 16'h120e, 16'h1221, 16'h1234, 16'h1247, 16'h125a, 16'h126d, 16'h1280, 16'h1293, 16'h12a6, 16'h12b9, 16'h12cc, 16'h12df, 16'h12f2, 16'h1305, 16'h1318, 16'h132b, 16'h133e, 16'h1351},
                                 {16'h1364, 16'h1377, 16'h138a, 16'h139d, 16'h13b0, 16'h13c3, 16'h13d6, 16'h13e9, 16'h13fc, 16'h140f, 16'h1422, 16'h1435, 16'h1448, 16'h145b, 16'h146e, 16'h1481, 16'h1494, 16'h14a7, 16'h14ba, 16'h14cd, 16'h14e0, 16'h14f3, 16'h1506, 16'h1519, 16'h152c, 16'h153f, 16'h1552, 16'h1565, 16'h1578, 16'h158b, 16'h159e, 16'h15b1, 16'h15c4, 16'h15d7, 16'h15ea, 16'h15fd, 16'h1610, 16'h1623, 16'h1636, 16'h1649, 16'h165c, 16'h166f, 16'h1682, 16'h1695, 16'h16a8, 16'h16bb, 16'h16ce, 16'h16e1, 16'h16f4, 16'h1707, 16'h171a, 16'h172d, 16'h1740, 16'h1753, 16'h1766, 16'h1779, 16'h178c, 16'h179f, 16'h17b2, 16'h17c5, 16'h17d8, 16'h17eb, 16'h17fe, 16'h1811},
                                 {16'h1824, 16'h1837, 16'h184a, 16'h185d, 16'h1870, 16'h1883, 16'h1896, 16'h18a9, 16'h18bc, 16'h18cf, 16'h18e2, 16'h18f5, 16'h1908, 16'h191b, 16'h192e, 16'h1941, 16'h1954, 16'h1967, 16'h197a, 16'h198d, 16'h19a0, 16'h19b3, 16'h19c6, 16'h19d9, 16'h19ec, 16'h19ff, 16'h1a12, 16'h1a25, 16'h1a38, 16'h1a4b, 16'h1a5e, 16'h1a71, 16'h1a84, 16'h1a97, 16'h1aaa, 16'h1abd, 16'h1ad0, 16'h1ae3, 16'h1af6, 16'h1b09, 16'h1b1c, 16'h1b2f, 16'h1b42, 16'h1b55, 16'h1b68, 16'h0d65, 16'h0d65, 16'h0d65, 16'h0d65, 16'h0d65, 16'h0d65, 16'h0d65, 16'h0d67, 16'h0d6b, 16'h0d6f, 16'h0d73, 16'h0d77, 16'h0d7b, 16'h0d7f, 16'h0d83, 16'h0d87, 16'h0d8b, 16'h0d8f, 16'h0d93},
                                 {16'h0d97, 16'h0d9b, 16'h0d9f, 16'h0da3, 16'h0da7, 16'h0dab, 16'h0daf, 16'h0db3, 16'h0db7, 16'h0dbb, 16'h0dbf, 16'h0dc3, 16'h0dc7, 16'h0dcb, 16'h0dcf, 16'h0dd3, 16'h0dd7, 16'h0ddb, 16'h0ddf, 16'h0de3, 16'h0de7, 16'h0deb, 16'h0def, 16'h0df3, 16'h0df7, 16'h0dfb, 16'h0dff, 16'h0e03, 16'h0e07, 16'h0e0b, 16'h0e0f, 16'h0e13, 16'h0e17, 16'h0e1b, 16'h0e1f, 16'h0e23, 16'h0e27, 16'h0e2b, 16'h0e2f, 16'h0e33, 16'h0e37, 16'h0e3b, 16'h0e3f, 16'h0e43, 16'h0e47, 16'h0e4b, 16'h0e4f, 16'h0e53, 16'h0e57, 16'h0e5b, 16'h0e5f, 16'h0e63, 16'h0e67, 16'h0e6b, 16'h0e6f, 16'h0e73, 16'h0e77, 16'h0e7b, 16'h0e7f, 16'h0e83, 16'h0e87, 16'h0e8b, 16'h0e8f, 16'h0e93},
                                 {16'h0e97, 16'h0e9b, 16'h0e9f, 16'h0ea3, 16'h0ea7, 16'h0eab, 16'h0eaf, 16'h0eb3, 16'h0eb7, 16'h0ebb, 16'h0ebf, 16'h0ec3, 16'h0ec7, 16'h0ecb, 16'h0ecf, 16'h0ed3, 16'h0ed7, 16'h0edb, 16'h0edf, 16'h0ee3, 16'h0ee7, 16'h0eeb, 16'h0eef, 16'h0ef3, 16'h0ef7, 16'h0efb, 16'h0eff, 16'h0f03, 16'h0f07, 16'h0f0b, 16'h0f0f, 16'h0f13, 16'h0f17, 16'h0f1b, 16'h0f1f, 16'h0f23, 16'h0f27, 16'h0f2b, 16'h0f2f, 16'h0f33, 16'h0f37, 16'h0f3b, 16'h0f3f, 16'h0f43, 16'h0f47, 16'h0f4b, 16'h0f4f, 16'h0f53, 16'h0f57, 16'h0f5b, 16'h0f5f, 16'h0f63, 16'h0f67, 16'h0f6b, 16'h0f6f, 16'h0f73, 16'h0f77, 16'h0f7b, 16'h0f7f, 16'h0f83, 16'h0f87, 16'h0f8b, 16'h0f8f, 16'h0f93},
                                 {16'h0f97, 16'h0f9b, 16'h0f9f, 16'h0fa3, 16'h0fa7, 16'h0fab, 16'h0faf, 16'h0fb3, 16'h0fb7, 16'h0fbb, 16'h0fbf, 16'h0fc3, 16'h0fc7, 16'h0fcb, 16'h0fcf, 16'h0fd3, 16'h0fd7, 16'h0fdb, 16'h0fdf, 16'h0fe3, 16'h0fe7, 16'h0feb, 16'h0fef, 16'h0ff3, 16'h0ff7, 16'h0ffb, 16'h0fff, 16'h1003, 16'h1007, 16'h100b, 16'h100f, 16'h1013, 16'h1017, 16'h101b, 16'h101f, 16'h1023, 16'h1027, 16'h102b, 16'h102f, 16'h1033, 16'h1037, 16'h103b, 16'h103f, 16'h1043, 16'h1047, 16'h104b, 16'h104f, 16'h1053, 16'h1057, 16'h105b, 16'h105f, 16'h1063, 16'h1067, 16'h106b, 16'h106f, 16'h1073, 16'h1077, 16'h107b, 16'h107f, 16'h1083, 16'h1087, 16'h108b, 16'h108f, 16'h1093},
                                 {16'h1097, 16'h109b, 16'h109f, 16'h10a3, 16'h10a7, 16'h10ab, 16'h10af, 16'h10b3, 16'h10b7, 16'h10bb, 16'h10bf, 16'h10c3, 16'h10c7, 16'h10cb, 16'h10cf, 16'h10d3, 16'h10d7, 16'h10db, 16'h10df, 16'h10e3, 16'h10e7, 16'h10eb, 16'h10ef, 16'h10f3, 16'h10f7, 16'h10fb, 16'h10ff, 16'h1103, 16'h1107, 16'h110b, 16'h110f, 16'h1113, 16'h1117, 16'h111b, 16'h111f, 16'h1123, 16'h10c6, 16'h10c4, 16'h10c2, 16'h10c0, 16'h10be, 16'h10bc, 16'h10ba, 16'h10b8, 16'h10b6, 16'h10b4, 16'h10b2, 16'h10b0, 16'h10ae, 16'h10ac, 16'h10aa, 16'h10a8, 16'h10a6, 16'h10a4, 16'h10a2, 16'h10a0, 16'h109e, 16'h109c, 16'h109a, 16'h1098, 16'h1096, 16'h1094, 16'h1092, 16'h1090},
                                 {16'h108e, 16'h108c, 16'h108a, 16'h1088, 16'h1086, 16'h1084, 16'h1082, 16'h1080, 16'h107e, 16'h107c, 16'h107a, 16'h1078, 16'h1076, 16'h1074, 16'h1072, 16'h1070, 16'h106e, 16'h106c, 16'h106a, 16'h1068, 16'h1066, 16'h1064, 16'h1062, 16'h1060, 16'h105e, 16'h105c, 16'h105a, 16'h1058, 16'h1056, 16'h1054, 16'h1052, 16'h1050, 16'h104e, 16'h104c, 16'h104a, 16'h1048, 16'h1046, 16'h1044, 16'h1042, 16'h1040, 16'h103e, 16'h103c, 16'h103a, 16'h1038, 16'h1036, 16'h1034, 16'h1032, 16'h1030, 16'h102e, 16'h102c, 16'h102a, 16'h1028, 16'h1026, 16'h1024, 16'h1022, 16'h1020, 16'h101e, 16'h101c, 16'h101a, 16'h1018, 16'h1016, 16'h1014, 16'h1012, 16'h1010},
                                 {16'h100e, 16'h100c, 16'h100a, 16'h1008, 16'h1006, 16'h1004, 16'h1002, 16'h1000, 16'h0ffe, 16'h0ffc, 16'h0ffa, 16'h0ff8, 16'h0ff6, 16'h0ff4, 16'h0ff2, 16'h0ff0, 16'h0fee, 16'h0fec, 16'h0fea, 16'h0fe8, 16'h0fe6, 16'h0fe4, 16'h0fe2, 16'h0fe0, 16'h0fde, 16'h0fdc, 16'h0fda, 16'h0fd8, 16'h0fd6, 16'h0fd4, 16'h0fd2, 16'h0fd0, 16'h0fce, 16'h0fcc, 16'h0fca, 16'h0fc8, 16'h0fc6, 16'h0fc4, 16'h0fc2, 16'h0fc0, 16'h0fbe, 16'h0fbc, 16'h0fba, 16'h0fb8, 16'h0fb6, 16'h0fb4, 16'h0fb2, 16'h0fb0, 16'h0fae, 16'h0fac, 16'h0faa, 16'h0fa8, 16'h0fa6, 16'h0fa4, 16'h0fa2, 16'h0fa0, 16'h0f9e, 16'h0f9c, 16'h0f9a, 16'h0f98, 16'h0f96, 16'h0f94, 16'h0f92, 16'h0f90},
                                 {16'h0f8e, 16'h0f8c, 16'h0f8a, 16'h0f88, 16'h0f86, 16'h0f84, 16'h0f82, 16'h0f80, 16'h0f7e, 16'h0f7c, 16'h0f7a, 16'h0f78, 16'h0f76, 16'h0f74, 16'h0f72, 16'h0f70, 16'h0f6e, 16'h0f6c, 16'h0f6a, 16'h0f68, 16'h0f66, 16'h0f64, 16'h0f62, 16'h0f60, 16'h0f5e, 16'h0f5c, 16'h0f5a, 16'h0f58, 16'h0f56, 16'h0f54, 16'h0f52, 16'h0f50, 16'h0f4e, 16'h0f4c, 16'h0f4a, 16'h0f48, 16'h0f46, 16'h0f44, 16'h0f42, 16'h0f40, 16'h0f3e, 16'h0f3c, 16'h0f3a, 16'h0f38, 16'h0f36, 16'h0f34, 16'h0f32, 16'h0f30, 16'h0f2e, 16'h0f2c, 16'h0f2a, 16'h0f28, 16'h0f26, 16'h0f24, 16'h0f22, 16'h0f20, 16'h0f1e, 16'h0f1c, 16'h0f1a, 16'h0f18, 16'h0f16, 16'h0f14, 16'h0f12, 16'h0f10},
                                 {16'h0f0e, 16'h0f0c, 16'h0f0a, 16'h0f08, 16'h0f06, 16'h0f04, 16'h0f02, 16'h0f00, 16'h0efe, 16'h0efc, 16'h0efa, 16'h0ef8, 16'h0ef6, 16'h0ef4, 16'h0ef2, 16'h0ef0, 16'h0eee, 16'h0eec, 16'h0eea, 16'h0ee8, 16'h0ee6, 16'h0ee4, 16'h0ee2, 16'h0ee0, 16'h0ede, 16'h0edc, 16'h0edc, 16'h0edc, 16'h0edc, 16'h0edc, 16'h0edc, 16'h0edc, 16'h0edc, 16'h0edc, 16'h0edc, 16'h0edc, 16'h0edc, 16'h0edc, 16'h0edc, 16'h0edc, 16'h0edc, 16'h0edc, 16'h0edc, 16'h0edc, 16'h0edc, 16'h0edc, 16'h0edc, 16'h0edc, 16'h0edc, 16'h0edc, 16'h0edc, 16'h0edc, 16'h0edc, 16'h0edf, 16'h0ee7, 16'h0eef, 16'h0ef7, 16'h0eff, 16'h0f07, 16'h0f0f, 16'h0f17, 16'h0f1f, 16'h0f27, 16'h0f2f},
                                 {16'h0f37, 16'h0f3f, 16'h0f47, 16'h0f4f, 16'h0f57, 16'h0f5f, 16'h0f67, 16'h0f6f, 16'h0f77, 16'h0f7f, 16'h0f87, 16'h0f8f, 16'h0f97, 16'h0f9f, 16'h0fa7, 16'h0faf, 16'h0fb7, 16'h0fbf, 16'h0fc7, 16'h0fcf, 16'h0fd7, 16'h0fdf, 16'h0fe7, 16'h0fef, 16'h0ff7, 16'h0fff, 16'h1007, 16'h100f, 16'h1017, 16'h101f, 16'h1027, 16'h102f, 16'h1037, 16'h103f, 16'h1047, 16'h104f, 16'h1057, 16'h105f, 16'h1067, 16'h106f, 16'h1077, 16'h107f, 16'h1087, 16'h108f, 16'h1097, 16'h109f, 16'h10a7, 16'h10af, 16'h10b7, 16'h10bf, 16'h10c7, 16'h10cf, 16'h10d7, 16'h10df, 16'h10e7, 16'h10ef, 16'h10f7, 16'h10ff, 16'h1107, 16'h110f, 16'h1117, 16'h111f, 16'h1127, 16'h112f},
                                 {16'h1137, 16'h113f, 16'h1147, 16'h114f, 16'h1157, 16'h115f, 16'h1167, 16'h116f, 16'h1177, 16'h117f, 16'h1187, 16'h118f, 16'h1197, 16'h119f, 16'h11a7, 16'h11af, 16'h11b7, 16'h11bf, 16'h11c7, 16'h11cf, 16'h11d7, 16'h11df, 16'h11e7, 16'h11ef, 16'h11f7, 16'h11ff, 16'h1207, 16'h120f, 16'h1217, 16'h121f, 16'h1227, 16'h122f, 16'h1237, 16'h123f, 16'h1247, 16'h124f, 16'h1257, 16'h125f, 16'h1267, 16'h126f, 16'h1277, 16'h127f, 16'h1287, 16'h128f, 16'h1297, 16'h129f, 16'h12a7, 16'h12af, 16'h12b7, 16'h12bf, 16'h12c7, 16'h12cf, 16'h12d7, 16'h12df, 16'h12e7, 16'h12ef, 16'h12f7, 16'h12ff, 16'h1307, 16'h130f, 16'h1317, 16'h131f, 16'h1327, 16'h132f},
                                 {16'h1337, 16'h133f, 16'h1347, 16'h134f, 16'h1357, 16'h135f, 16'h1367, 16'h136f, 16'h1377, 16'h137f, 16'h1387, 16'h138f, 16'h1397, 16'h139f, 16'h13a7, 16'h13af, 16'h13b7, 16'h13bf, 16'h13c7, 16'h13cf, 16'h13d7, 16'h13df, 16'h13e7, 16'h13ef, 16'h13f7, 16'h13ff, 16'h1407, 16'h140f, 16'h1417, 16'h141f, 16'h1427, 16'h142f, 16'h1437, 16'h143f, 16'h1447, 16'h144f, 16'h1457, 16'h145f, 16'h1467, 16'h146f, 16'h1477, 16'h147f, 16'h1487, 16'h148f, 16'h1497, 16'h149f, 16'h14a7, 16'h14af, 16'h14b7, 16'h14bf, 16'h14c7, 16'h14cf, 16'h14d7, 16'h14df, 16'h14e7, 16'h14ef, 16'h14f7, 16'h14ff, 16'h1507, 16'h150f, 16'h1517, 16'h151f, 16'h1527, 16'h152f},
                                 {16'h1537, 16'h153f, 16'h1547, 16'h154f, 16'h1557, 16'h155f, 16'h1567, 16'h156f, 16'h1577, 16'h157f, 16'h1587, 16'h158f, 16'h1597, 16'h159f, 16'h15a7, 16'h15af, 16'h15b7, 16'h15bf, 16'h15c7, 16'h15cf, 16'h15d7, 16'h15df, 16'h15e7, 16'h15ef, 16'h15f7, 16'h15ff, 16'h1607, 16'h160f, 16'h1617, 16'h161f, 16'h1627, 16'h162f, 16'h1637, 16'h163f, 16'h1647, 16'h164f, 16'h1657, 16'h165f, 16'h1667, 16'h166f, 16'h1677, 16'h167f, 16'h1687, 16'h168f, 16'h1697, 16'h169f, 16'h16a7, 16'h16af, 16'h16b7, 16'h16bf, 16'h16c7, 16'h16cf, 16'h16d7, 16'h16df, 16'h16e7, 16'h16ef, 16'h16f7, 16'h16ff, 16'h1707, 16'h170f, 16'h1717, 16'h171f, 16'h1727, 16'h172f},
                                 {16'h1737, 16'h173f, 16'h1747, 16'h174f, 16'h1757, 16'h175f, 16'h1767, 16'h176f, 16'h1777, 16'h177f, 16'h1787, 16'h178f, 16'h1797, 16'h179f, 16'h17a7, 16'h17af, 16'h17b7, 16'h17bf, 16'h17c7, 16'h17cf, 16'h17d7, 16'h17df, 16'h17e7, 16'h17ef, 16'h17f7, 16'h17ff, 16'h1807, 16'h180f, 16'h1817, 16'h181f, 16'h1827, 16'h182f, 16'h1837, 16'h183f, 16'h1847, 16'h184f, 16'h1857, 16'h185f, 16'h1867, 16'h186f, 16'h1877, 16'h187f, 16'h1887, 16'h188f, 16'h1897, 16'h189f, 16'h18a7, 16'h18af, 16'h18b7, 16'h18bf, 16'h18c7, 16'h18cf, 16'h18d7, 16'h18df, 16'h18e7, 16'h18ef, 16'h18f7, 16'h18ff, 16'h1907, 16'h190f, 16'h1917, 16'h191f, 16'h1927, 16'h192f},
                                 {16'h1937, 16'h193f, 16'h1947, 16'h194f, 16'h1957, 16'h195f, 16'h1967, 16'h196f, 16'h1977, 16'h197f, 16'h1987, 16'h198f, 16'h1997, 16'h199f, 16'h19a7, 16'h19af, 16'h19b7, 16'h19bf, 16'h19c7, 16'h19cf, 16'h19d7, 16'h19df, 16'h19e7, 16'h19ef, 16'h19f7, 16'h19ff, 16'h1a07, 16'h1a0f, 16'h1a17, 16'h1a1f, 16'h1a27, 16'h1a2f, 16'h1a37, 16'h1a3f, 16'h1a47, 16'h1a4f, 16'h1a57, 16'h1a5f, 16'h1a67, 16'h1a6f, 16'h1a77, 16'h1a7f, 16'h1a87, 16'h1a8f, 16'h1a97, 16'h1a9f, 16'h1aa7, 16'h1aaf, 16'h1ab7, 16'h1abf, 16'h1ac7, 16'h1acf, 16'h1ad7, 16'h1adf, 16'h1ae7, 16'h1aef, 16'h1af7, 16'h1aff, 16'h1b07, 16'h1b0f, 16'h1b17, 16'h1b1f, 16'h1b27, 16'h1b2f},
                                 {16'h1b37, 16'h1b3f, 16'h1b47, 16'h1b4f, 16'h1b57, 16'h1b5f, 16'h1b67, 16'h1b6f, 16'h1b77, 16'h1b7f, 16'h1b87, 16'h1b8f, 16'h1b97, 16'h1b9f, 16'h1ba7, 16'h1baf, 16'h1bb7, 16'h1bbf, 16'h1bc7, 16'h1bcf, 16'h1bd7, 16'h1bdf, 16'h1be7, 16'h1bef, 16'h1bf7, 16'h1bff, 16'h1c07, 16'h1c0f, 16'h1c17, 16'h1c1f, 16'h1c27, 16'h1c2f, 16'h1c37, 16'h1c3f, 16'h1c47, 16'h1c4f, 16'h1c57, 16'h1c5f, 16'h1c67, 16'h1c6f, 16'h1c77, 16'h1c7f, 16'h1c87, 16'h1c8f, 16'h1c97, 16'h1c9f, 16'h1ca7, 16'h1caf, 16'h1cb7, 16'h1cbf, 16'h1cc7, 16'h1ccf, 16'h1cd7, 16'h1cdf, 16'h1ce7, 16'h1cef, 16'h1cf7, 16'h1cff, 16'h1d07, 16'h1d0f, 16'h1d17, 16'h1d1f, 16'h1d27, 16'h1d2f},
                                 {16'h1d37, 16'h1d3f, 16'h1d47, 16'h1d4f, 16'h1d57, 16'h1d5f, 16'h1d67, 16'h1d6f, 16'h1d77, 16'h1d7f, 16'h1d87, 16'h1d8f, 16'h1d97, 16'h1d9f, 16'h1da7, 16'h1daf, 16'h1db7, 16'h1dbf, 16'h1dc7, 16'h1dcf, 16'h1dd7, 16'h1ddf, 16'h1de7, 16'h1def, 16'h1df7, 16'h1dff, 16'h1e07, 16'h1e0f, 16'h1e17, 16'h1e1f, 16'h1e27, 16'h1e2f, 16'h1e37, 16'h1e3f, 16'h1e47, 16'h1e4f, 16'h1e57, 16'h1e5f, 16'h1e67, 16'h1e6f, 16'h1e77, 16'h1e7f, 16'h1e87, 16'h1e8f, 16'h1e97, 16'h1e9f, 16'h1ea7, 16'h1eaf, 16'h1eb7, 16'h1ebf, 16'h1ec7, 16'h1ecf, 16'h1ed7, 16'h1edf, 16'h1ee7, 16'h1eef, 16'h1ef7, 16'h1eff, 16'h1f07, 16'h1f0f, 16'h1f17, 16'h1f1f, 16'h1f27, 16'h1f2f},
                                 {16'h1f37, 16'h1f3f, 16'h1f47, 16'h1f4f, 16'h1f57, 16'h1f57, 16'h1f3d, 16'h1f10, 16'h1ee3, 16'h1eb6, 16'h1e89, 16'h1e5c, 16'h1e2f, 16'h1e02, 16'h1dd5, 16'h1da8, 16'h1d7b, 16'h1d4e, 16'h1d21, 16'h1cf4, 16'h1cc7, 16'h1c9a, 16'h1c6d, 16'h1c40, 16'h1c13, 16'h1be6, 16'h1bb9, 16'h1b8c, 16'h1b5f, 16'h1b32, 16'h1b05, 16'h1ad8, 16'h1aab, 16'h1a7e, 16'h1a51, 16'h1a24, 16'h19f7, 16'h19ca, 16'h199d, 16'h1970, 16'h1943, 16'h1916, 16'h18e9, 16'h18bc, 16'h188f, 16'h1862, 16'h1835, 16'h1808, 16'h17db, 16'h17ae, 16'h1781, 16'h1754, 16'h1727, 16'h16fa, 16'h16cd, 16'h16a0, 16'h1673, 16'h1646, 16'h1619, 16'h15ec, 16'h15bf, 16'h1592, 16'h1565, 16'h1538},
                                 {16'h150b, 16'h14de, 16'h14b1, 16'h1484, 16'h1457, 16'h142a, 16'h13fd, 16'h13d0, 16'h13a3, 16'h1376, 16'h1349, 16'h131c, 16'h12ef, 16'h12c2, 16'h1295, 16'h1268, 16'h123b, 16'h120e, 16'h11e1, 16'h11b4, 16'h1187, 16'h115a, 16'h112d, 16'h1100, 16'h10d3, 16'h10a6, 16'h1079, 16'h104c, 16'h101f, 16'h0ff2, 16'h0fc5, 16'h0f98, 16'h0f6b, 16'h0f3e, 16'h0f11, 16'h0ee4, 16'h0eb7, 16'h0e8a, 16'h0e5d, 16'h0e30, 16'h0e03, 16'h0dd6, 16'h0da9, 16'h0d7c, 16'h0d4f, 16'h0d22, 16'h0cf5, 16'h0cc8, 16'h0c9b, 16'h0c6e, 16'h0c41, 16'h0c14, 16'h0be7, 16'h0bba, 16'h0b8d, 16'h0b60, 16'h0b33, 16'h0b06, 16'h0ad9, 16'h0aac, 16'h0a7f, 16'h0a52, 16'h0a25, 16'h09f8},
                                 {16'h09cb, 16'h099e, 16'h0971, 16'h0944, 16'h0917, 16'h08ea, 16'h08bd, 16'h0890, 16'h0863, 16'h0836, 16'h0809, 16'h07dc, 16'h07af, 16'h0782, 16'h0755, 16'h0728, 16'h06fb, 16'h06ce, 16'h06a1, 16'h0674, 16'h2764, 16'h2717, 16'h26f5, 16'h26d3, 16'h26b1, 16'h268f, 16'h266d, 16'h264b, 16'h2629, 16'h2607, 16'h25e5, 16'h25c3, 16'h25a1, 16'h257f, 16'h255d, 16'h253b, 16'h2519, 16'h24f7, 16'h24d5, 16'h24b3, 16'h2491, 16'h246f, 16'h244d, 16'h242b, 16'h2409, 16'h23e7, 16'h23c5, 16'h23a3, 16'h2381, 16'h235f, 16'h233d, 16'h231b, 16'h22f9, 16'h22d7, 16'h22b5, 16'h2293, 16'h2271, 16'h224f, 16'h222d, 16'h220b, 16'h21e9, 16'h21c7, 16'h21a5, 16'h2183},
                                 {16'h2161, 16'h213f, 16'h211d, 16'h20fb, 16'h20d9, 16'h20b7, 16'h2095, 16'h2073, 16'h2051, 16'h202f, 16'h200d, 16'h1feb, 16'h1fc9, 16'h1fa7, 16'h1f85, 16'h1f63, 16'h1f41, 16'h1f1f, 16'h1efd, 16'h1edb, 16'h1eb9, 16'h1e97, 16'h1e75, 16'h1e53, 16'h1e31, 16'h1e0f, 16'h1ded, 16'h1dcb, 16'h1da9, 16'h1d87, 16'h1d65, 16'h1d43, 16'h1d21, 16'h1cff, 16'h1cdd, 16'h1cbb, 16'h1c99, 16'h1c77, 16'h1c55, 16'h1c33, 16'h1c11, 16'h1bef, 16'h1bcd, 16'h1bab, 16'h1b89, 16'h1b67, 16'h1b45, 16'h1b23, 16'h1b01, 16'h1adf, 16'h1abd, 16'h1a9b, 16'h1a79, 16'h1a57, 16'h1a35, 16'h1a13, 16'h19f1, 16'h19cf, 16'h19ad, 16'h198b, 16'h1969, 16'h1947, 16'h1925, 16'h1903},
                                 {16'h18e1, 16'h18bf, 16'h189d, 16'h187b, 16'h1859, 16'h1837, 16'h1815, 16'h17f3, 16'h17d1, 16'h17af, 16'h178d, 16'h176b, 16'h1749, 16'h1727, 16'h1705, 16'h16e3, 16'h16c1, 16'h169f, 16'h167d, 16'h165b, 16'h1639, 16'h1617, 16'h15f5, 16'h15d3, 16'h15b1, 16'h158f, 16'h156d, 16'h154b, 16'h1529, 16'h1507, 16'h14e5, 16'h14c3, 16'h14a1, 16'h147f, 16'h145d, 16'h143b, 16'h1419, 16'h13f7, 16'h13d5, 16'h13b3, 16'h1391, 16'h136f, 16'h134d, 16'h132b, 16'h1309, 16'h12e7, 16'h12c5, 16'h12a3, 16'h1281, 16'h125f, 16'h123d, 16'h121b, 16'h11f9, 16'h11d7, 16'h11b5, 16'h1193, 16'h1171, 16'h114f, 16'h112d, 16'h110b, 16'h10e9, 16'h10c7, 16'h10a5, 16'h1083},
                                 {16'h1061, 16'h103f, 16'h101d, 16'h0ffb, 16'h0fd9, 16'h0fb7, 16'h0f95, 16'h0f73, 16'h0f51, 16'h0f2f, 16'h0f0d, 16'h0eeb, 16'h0ec9, 16'h0ea7, 16'h0e85, 16'h0e63, 16'h0e41, 16'h0e1f, 16'h0dfd, 16'h0ddb, 16'h0db9, 16'h0d97, 16'h0d75, 16'h0d53, 16'h0d31, 16'h0d0f, 16'h0ced, 16'h0ccb, 16'h0ca9, 16'h0d1a, 16'h0d56, 16'h0d92, 16'h0dce, 16'h0e0a, 16'h0e46, 16'h0e82, 16'h0ebe, 16'h0efa, 16'h0f36, 16'h0f72, 16'h0fae, 16'h0fea, 16'h1026, 16'h1062, 16'h109e, 16'h10da, 16'h1116, 16'h1152, 16'h118e, 16'h11ca, 16'h1206, 16'h1242, 16'h127e, 16'h12ba, 16'h12f6, 16'h1332, 16'h136e, 16'h13aa, 16'h13e6, 16'h1422, 16'h145e, 16'h149a, 16'h14d6, 16'h1512},
                                 {16'h154e, 16'h158a, 16'h15c6, 16'h1602, 16'h163e, 16'h167a, 16'h16b6, 16'h16f2, 16'h172e, 16'h176a, 16'h17a6, 16'h17e2, 16'h181e, 16'h185a, 16'h1896, 16'h18d2, 16'h190e, 16'h194a, 16'h1986, 16'h19c2, 16'h19fe, 16'h1a3a, 16'h1a76, 16'h1ab2, 16'h1aee, 16'h1b2a, 16'h1b66, 16'h1ba2, 16'h1bde, 16'h1c1a, 16'h1c56, 16'h1c92, 16'h1cce, 16'h1d0a, 16'h1d46, 16'h1d82, 16'h1dbe, 16'h1dfa, 16'h1e36, 16'h1e72, 16'h1eae, 16'h1eea, 16'h1f26, 16'h1f62, 16'h1f9e, 16'h1fda, 16'h2016, 16'h2052, 16'h208e, 16'h20ca, 16'h2106, 16'h2142, 16'h217e, 16'h21ba, 16'h21f6, 16'h2232, 16'h226e, 16'h22aa, 16'h22e6, 16'h2322, 16'h235e, 16'h239a, 16'h23d6, 16'h2412},
                                 {16'h244e, 16'h248a, 16'h24c6, 16'h2502, 16'h253e, 16'h257a, 16'h25b6, 16'h25f2, 16'h262e, 16'h266a, 16'h26a6, 16'h26e2, 16'h271e, 16'h275a, 16'h2796, 16'h27d2, 16'h280e, 16'h284a, 16'h2886, 16'h28c2, 16'h28fe, 16'h293a, 16'h2976, 16'h29b2, 16'h29ee, 16'h2a2a, 16'h2a66, 16'h2aa2, 16'h2ade, 16'h2b1a, 16'h2b56, 16'h2b92, 16'h2bce, 16'h2c0a, 16'h2c46, 16'h2c82, 16'h2cbe, 16'h2cfa, 16'h2d36, 16'h2d72, 16'h2dae, 16'h2dea, 16'h2e26, 16'h2e62, 16'h2e9e, 16'h2eda, 16'h2f16, 16'h2f52, 16'h2f8e, 16'h2fca, 16'h3006, 16'h3042, 16'h307e, 16'h30ba, 16'h30f6, 16'h3132, 16'h316e, 16'h31aa, 16'h31e6, 16'h3222, 16'h325e, 16'h329a, 16'h32d6, 16'h3312},
                                 {16'h334e, 16'h338a, 16'h33c6, 16'h3402, 16'h343e, 16'h347a, 16'h34b6, 16'h34f2, 16'h352e, 16'h356a, 16'h35a6, 16'h35e2, 16'h361e, 16'h365a, 16'h3696, 16'h36d2, 16'h370e, 16'h374a, 16'h3786, 16'h37c2, 16'h37fe, 16'h383a, 16'h3876, 16'h38b2, 16'h38ee, 16'h392a, 16'h3966, 16'h39a2, 16'h39de, 16'h3a1a, 16'h3a56, 16'h3a92, 16'h3ace, 16'h3b0a, 16'h3b46, 16'h3b82, 16'h3bbe, 16'h3bfa, 16'h3c36, 16'h3c72, 16'h3cae, 16'h3cea, 16'h3c73, 16'h3c69, 16'h3c5f, 16'h3c55, 16'h3c4b, 16'h3c41, 16'h3c37, 16'h3c2d, 16'h3c23, 16'h3c19, 16'h3c0f, 16'h3c05, 16'h3bfb, 16'h3bf1, 16'h3be7, 16'h3bdd, 16'h3bd3, 16'h3bc9, 16'h3bbf, 16'h3bb5, 16'h3bab, 16'h3ba1},
                                 {16'h3b97, 16'h3b8d, 16'h3b83, 16'h3b79, 16'h3b6f, 16'h3b65, 16'h3b5b, 16'h3b51, 16'h3b47, 16'h3b3d, 16'h3b33, 16'h3b29, 16'h3b1f, 16'h3b15, 16'h3b0b, 16'h3b01, 16'h3af7, 16'h3aed, 16'h3ae3, 16'h3ad9, 16'h3acf, 16'h3ac5, 16'h3abb, 16'h3ab1, 16'h3aa7, 16'h3a9d, 16'h3a93, 16'h3a89, 16'h3a7f, 16'h3a75, 16'h3a6b, 16'h3a61, 16'h3a57, 16'h3a4d, 16'h3a43, 16'h3a39, 16'h3a2f, 16'h3a25, 16'h3a1b, 16'h3a11, 16'h3a07, 16'h39fd, 16'h39f3, 16'h39e9, 16'h39df, 16'h39d5, 16'h39cb, 16'h39c1, 16'h39b7, 16'h39ad, 16'h39a3, 16'h3999, 16'h398f, 16'h3985, 16'h397b, 16'h3971, 16'h3967, 16'h395d, 16'h3953, 16'h3949, 16'h393f, 16'h3935, 16'h392b, 16'h3921},
                                 {16'h3917, 16'h390d, 16'h3903, 16'h38f9, 16'h38ef, 16'h38e5, 16'h38db, 16'h38d1, 16'h38c7, 16'h38bd, 16'h38b3, 16'h38a9, 16'h389f, 16'h3895, 16'h388b, 16'h3881, 16'h3877, 16'h386d, 16'h3863, 16'h3859, 16'h384f, 16'h3845, 16'h383b, 16'h3831, 16'h3827, 16'h381d, 16'h3813, 16'h3809, 16'h37ff, 16'h37f5, 16'h37eb, 16'h37e1, 16'h37d7, 16'h37cd, 16'h37c3, 16'h37b9, 16'h37af, 16'h37a5, 16'h379b, 16'h3791, 16'h3787, 16'h377d, 16'h3773, 16'h3769, 16'h375f, 16'h3755, 16'h374b, 16'h3741, 16'h3737, 16'h372d, 16'h3723, 16'h3719, 16'h370f, 16'h3705, 16'h36fb, 16'h36f1, 16'h36e7, 16'h36dd, 16'h36d3, 16'h36c9, 16'h36bf, 16'h36b5, 16'h36ab, 16'h36a1},
                                 {16'h3697, 16'h368d, 16'h3683, 16'h3679, 16'h366f, 16'h3665, 16'h365b, 16'h3651, 16'h3647, 16'h363d, 16'h3633, 16'h3629, 16'h361f, 16'h3615, 16'h360b, 16'h3601, 16'h35f7, 16'h35ed, 16'h35e3, 16'h35d9, 16'h35cf, 16'h35c5, 16'h35bb, 16'h35b1, 16'h35a7, 16'h359d, 16'h3593, 16'h3589, 16'h357f, 16'h3575, 16'h356b, 16'h3561, 16'h3557, 16'h354d, 16'h3543, 16'h3539, 16'h352f, 16'h3525, 16'h351b, 16'h3511, 16'h3507, 16'h34fd, 16'h34f3, 16'h34e9, 16'h34df, 16'h34d5, 16'h34cb, 16'h34c1, 16'h34b7, 16'h34ad, 16'h34a3, 16'h3499, 16'h348f, 16'h3485, 16'h347b, 16'h3471, 16'h3467, 16'h345d, 16'h3453, 16'h3449, 16'h343f, 16'h3435, 16'h342b, 16'h3421},
                                 {16'h3417, 16'h340d, 16'h3403, 16'h33f9, 16'h33ef, 16'h33e5, 16'h33db, 16'h33d1, 16'h33c7, 16'h33bd, 16'h33b3, 16'h33a9, 16'h339f, 16'h3395, 16'h338b, 16'h3381, 16'h3377, 16'h336d, 16'h3363, 16'h3359, 16'h334f, 16'h3345, 16'h333b, 16'h3331, 16'h3327, 16'h331d, 16'h3313, 16'h3309, 16'h32ff, 16'h32f5, 16'h32eb, 16'h32e1, 16'h32d7, 16'h32cd, 16'h32c3, 16'h32b9, 16'h32af, 16'h32a5, 16'h329b, 16'h3291, 16'h3287, 16'h327d, 16'h3273, 16'h3269, 16'h325f, 16'h3255, 16'h324b, 16'h3241, 16'h3237, 16'h322d, 16'h3223, 16'h3219, 16'h320f, 16'h3205, 16'h31fb, 16'h31f1, 16'h31e7, 16'h31dd, 16'h31d3, 16'h31c9, 16'h31bf, 16'h31b5, 16'h31ab, 16'h31a1},
                                 {16'h3197, 16'h318d, 16'h3183, 16'h3179, 16'h316f, 16'h3165, 16'h315b, 16'h3151, 16'h3147, 16'h313d, 16'h3133, 16'h3129, 16'h311f, 16'h3115, 16'h310b, 16'h3101, 16'h30f7, 16'h30ed, 16'h30e3, 16'h30d9, 16'h30cf, 16'h30c5, 16'h30bb, 16'h30b1, 16'h30a7, 16'h309d, 16'h3093, 16'h3089, 16'h307f, 16'h3075, 16'h306b, 16'h3061, 16'h3057, 16'h304d, 16'h3043, 16'h3039, 16'h302f, 16'h3025, 16'h301b, 16'h3011, 16'h3007, 16'h2ffd, 16'h2ff3, 16'h2fe9, 16'h2fdf, 16'h2fd5, 16'h2fcb, 16'h2fc1, 16'h2fb7, 16'h2fad, 16'h2fa3, 16'h2f99, 16'h2f8f, 16'h2f85, 16'h2f7b, 16'h2f71, 16'h2f67, 16'h2f5d, 16'h2f53, 16'h2f49, 16'h2f3f, 16'h2f35, 16'h2f2b, 16'h2f21},
                                 {16'h2f17, 16'h2f0d, 16'h2f03, 16'h2ef9, 16'h2eef, 16'h2ee5, 16'h2edb, 16'h2ed1, 16'h2ec7, 16'h2ebd, 16'h2eb3, 16'h2ea9, 16'h2e9f, 16'h2e95, 16'h2e8b, 16'h2e81, 16'h2e77, 16'h2e6d, 16'h2e63, 16'h2e59, 16'h2e4f, 16'h2e45, 16'h2e3b, 16'h2e31, 16'h2e27, 16'h2e1d, 16'h2e13, 16'h2e09, 16'h2dff, 16'h2df5, 16'h2deb, 16'h2de1, 16'h2dd7, 16'h2dcd, 16'h2dc3, 16'h2db9, 16'h2daf, 16'h2da5, 16'h2d9b, 16'h2d91, 16'h2d87, 16'h2d7d, 16'h2d73, 16'h2d69, 16'h2d5f, 16'h2d55, 16'h2d4b, 16'h2d41, 16'h2d37, 16'h2d2d, 16'h2d23, 16'h2d19, 16'h2d0f, 16'h2d05, 16'h2cfb, 16'h2cf1, 16'h2ce7, 16'h2cdd, 16'h2cd3, 16'h2cc9, 16'h2cbf, 16'h2cb5, 16'h2cab, 16'h2ca1},
                                 {16'h2c97, 16'h2c8d, 16'h2c83, 16'h2c79, 16'h2c6f, 16'h2c65, 16'h2c5b, 16'h2c51, 16'h2c47, 16'h2c3d, 16'h2c33, 16'h2c29, 16'h2c1f, 16'h2c15, 16'h2c0b, 16'h2c01, 16'h2bf7, 16'h2bed, 16'h2be3, 16'h2bd9, 16'h2bcf, 16'h2bc5, 16'h2bbb, 16'h2bb1, 16'h2ba7, 16'h2b9d, 16'h2b93, 16'h2b89, 16'h2b7f, 16'h2b75, 16'h2b6b, 16'h2b61, 16'h2b57, 16'h2b4d, 16'h2b43, 16'h2b39, 16'h2b2f, 16'h2b25, 16'h2b1b, 16'h2b11, 16'h2b07, 16'h2afd, 16'h2af3, 16'h2ae9, 16'h2adf, 16'h2ad5, 16'h2acb, 16'h2ac1, 16'h2ab7, 16'h2aad, 16'h2aa3, 16'h2a99, 16'h2a8f, 16'h2a85, 16'h2a7b, 16'h2a71, 16'h2a67, 16'h2a5d, 16'h2a53, 16'h2a49, 16'h2a3f, 16'h2a35, 16'h2a2b, 16'h2a21},
                                 {16'h2a17, 16'h2a0d, 16'h2a03, 16'h29f9, 16'h29ef, 16'h29e5, 16'h29db, 16'h29d1, 16'h29c7, 16'h29bd, 16'h29b3, 16'h29a9, 16'h299f, 16'h2995, 16'h298b, 16'h2981, 16'h2977, 16'h296d, 16'h2963, 16'h2959, 16'h294f, 16'h2945, 16'h293b, 16'h2931, 16'h2927, 16'h291d, 16'h2913, 16'h2909, 16'h28ff, 16'h28f5, 16'h28eb, 16'h28e1, 16'h28d7, 16'h28cd, 16'h28c3, 16'h28b9, 16'h28af, 16'h28a5, 16'h289b, 16'h2891, 16'h2887, 16'h287d, 16'h2873, 16'h2869, 16'h285f, 16'h2855, 16'h284b, 16'h2841, 16'h2837, 16'h282d, 16'h2823, 16'h2819, 16'h280f, 16'h2805, 16'h27fb, 16'h27f1, 16'h27e7, 16'h27dd, 16'h27d3, 16'h27c9, 16'h27bf, 16'h27b5, 16'h27ab, 16'h27a1},
                                 {16'h2797, 16'h278d, 16'h2783, 16'h2779, 16'h276f, 16'h2765, 16'h275b, 16'h2731, 16'h26fc, 16'h26c7, 16'h2692, 16'h265d, 16'h2628, 16'h25f3, 16'h25be, 16'h2589, 16'h2554, 16'h251f, 16'h24ea, 16'h24b5, 16'h2480, 16'h244b, 16'h2416, 16'h23e1, 16'h23ac, 16'h2377, 16'h2342, 16'h230d, 16'h22d8, 16'h22a3, 16'h226e, 16'h2239, 16'h2204, 16'h21cf, 16'h219a, 16'h2165, 16'h2130, 16'h20fb, 16'h20c6, 16'h2091, 16'h205c, 16'h2027, 16'h1ff2, 16'h1fbd, 16'h1f88, 16'h1f53, 16'h1f1e, 16'h1ee9, 16'h1eb4, 16'h1e7f, 16'h1e7f, 16'h1e7f, 16'h1e7f, 16'h1e7f, 16'h1e7f, 16'h1e76, 16'h1e65, 16'h1e54, 16'h1e43, 16'h1e32, 16'h1e21, 16'h1e10, 16'h1dff, 16'h1dee},
                                 {16'h1ddd, 16'h1dcc, 16'h1dbb, 16'h1daa, 16'h1d99, 16'h1d88, 16'h1d77, 16'h1d66, 16'h1d55, 16'h1d44, 16'h1d33, 16'h1d22, 16'h1d11, 16'h1d00, 16'h1cef, 16'h1cde, 16'h1ccd, 16'h1cbc, 16'h1cab, 16'h1c9a, 16'h1c89, 16'h1c78, 16'h1c67, 16'h1c56, 16'h1c45, 16'h1c34, 16'h1c23, 16'h1c12, 16'h1c01, 16'h1bf0, 16'h1bdf, 16'h1bce, 16'h1bbd, 16'h1bac, 16'h1b9b, 16'h1b8a, 16'h1b79, 16'h1b68, 16'h1b57, 16'h1b46, 16'h1b35, 16'h1b24, 16'h1b13, 16'h1b02, 16'h1af1, 16'h1ae0, 16'h1acf, 16'h1abe, 16'h1aad, 16'h1a9c, 16'h1a8b, 16'h1a7a, 16'h1a69, 16'h1a58, 16'h1a47, 16'h1a36, 16'h1a25, 16'h1a14, 16'h1a03, 16'h19f2, 16'h19e1, 16'h19d0, 16'h19bf, 16'h19ae},
                                 {16'h199d, 16'h198c, 16'h197b, 16'h196a, 16'h1959, 16'h1948, 16'h1937, 16'h1926, 16'h1915, 16'h1904, 16'h18f3, 16'h18e2, 16'h18d1, 16'h18c0, 16'h18af, 16'h189e, 16'h188d, 16'h187c, 16'h186b, 16'h185a, 16'h1849, 16'h1838, 16'h1827, 16'h1816, 16'h1805, 16'h17f4, 16'h17e3, 16'h17d2, 16'h17c1, 16'h17b0, 16'h179f, 16'h178e, 16'h177d, 16'h176c, 16'h175b, 16'h174a, 16'h1739, 16'h1728, 16'h1717, 16'h1706, 16'h16f5, 16'h16e4, 16'h16d3, 16'h16c2, 16'h16b1, 16'h16a0, 16'h168f, 16'h167e, 16'h166d, 16'h165c, 16'h164b, 16'h163a, 16'h1629, 16'h1618, 16'h1607, 16'h15f6, 16'h15e5, 16'h15d4, 16'h15c3, 16'h15b2, 16'h15a1, 16'h1590, 16'h157f, 16'h156e},
                                 {16'h155d, 16'h154c, 16'h153b, 16'h152a, 16'h1519, 16'h1508, 16'h14f7, 16'h14e6, 16'h14d5, 16'h14c4, 16'h14b3, 16'h14a2, 16'h1491, 16'h1480, 16'h146f, 16'h145e, 16'h144d, 16'h143c, 16'h142b, 16'h141a, 16'h1409, 16'h13f8, 16'h13e7, 16'h13d6, 16'h13c5, 16'h13b4, 16'h13a3, 16'h1392, 16'h1381, 16'h1370, 16'h135f, 16'h134e, 16'h133d, 16'h132c, 16'h131b, 16'h130a, 16'h12f9, 16'h12e8, 16'h12d7, 16'h12c6, 16'h12b5, 16'h12a4, 16'h1293, 16'h1282, 16'h1271, 16'h1260, 16'h124f, 16'h123e, 16'h122d, 16'h121c, 16'h120b, 16'h11fa, 16'h11e9, 16'h11d8, 16'h11c7, 16'h11b6, 16'h11a5, 16'h1194, 16'h1183, 16'h1172, 16'h1161, 16'h1150, 16'h113f, 16'h112e},
                                 {16'h111d, 16'h110c, 16'h10fb, 16'h10ea, 16'h10d9, 16'h10c8, 16'h10b7, 16'h10a6, 16'h1095, 16'h1084, 16'h1073, 16'h1062, 16'h1051, 16'h1040, 16'h102f, 16'h101e, 16'h100d, 16'h0ffc, 16'h0feb, 16'h0fda, 16'h0fc9, 16'h0fb8, 16'h0fa7, 16'h0f96, 16'h0f85, 16'h0f74, 16'h0f63, 16'h0f52, 16'h0f41, 16'h0f30, 16'h0f1f, 16'h0f0e, 16'h0efd, 16'h0eec, 16'h0edb, 16'h0edb, 16'h0edb, 16'h0edb, 16'h0edb, 16'h0edb, 16'h0eec, 16'h0f08, 16'h0f24, 16'h0f40, 16'h0f5c, 16'h0f78, 16'h0f94, 16'h0fb0, 16'h0fcc, 16'h0fe8, 16'h1004, 16'h1020, 16'h103c, 16'h1058, 16'h1074, 16'h1090, 16'h10ac, 16'h10c8, 16'h10e4, 16'h1100, 16'h111c, 16'h1138, 16'h1154, 16'h1170},
                                 {16'h118c, 16'h11a8, 16'h11c4, 16'h11e0, 16'h11fc, 16'h1218, 16'h1234, 16'h1250, 16'h126c, 16'h1288, 16'h12a4, 16'h12c0, 16'h12dc, 16'h12f8, 16'h1314, 16'h1330, 16'h134c, 16'h1368, 16'h1384, 16'h13a0, 16'h13bc, 16'h13d8, 16'h13f4, 16'h1410, 16'h142c, 16'h1448, 16'h1464, 16'h1480, 16'h149c, 16'h14b8, 16'h14d4, 16'h14f0, 16'h150c, 16'h1528, 16'h1544, 16'h1560, 16'h157c, 16'h1598, 16'h15b4, 16'h15d0, 16'h15ec, 16'h1608, 16'h1624, 16'h1640, 16'h165c, 16'h1678, 16'h1694, 16'h16b0, 16'h16cc, 16'h16e8, 16'h1704, 16'h1720, 16'h173c, 16'h1758, 16'h1774, 16'h1790, 16'h17ac, 16'h17c8, 16'h17e4, 16'h1800, 16'h181c, 16'h1838, 16'h1854, 16'h1870},
                                 {16'h188c, 16'h18a8, 16'h18c4, 16'h18e0, 16'h18fc, 16'h1918, 16'h1934, 16'h1950, 16'h196c, 16'h1988, 16'h19a4, 16'h19c0, 16'h19dc, 16'h19f8, 16'h1a14, 16'h1a30, 16'h1a4c, 16'h1a68, 16'h1a84, 16'h1aa0, 16'h1abc, 16'h1ad8, 16'h1af4, 16'h1b10, 16'h1b2c, 16'h1b48, 16'h1b64, 16'h1b80, 16'h1b9c, 16'h1bb8, 16'h1bd4, 16'h1bf0, 16'h1c0c, 16'h1c28, 16'h1c44, 16'h1c60, 16'h1c7c, 16'h1c98, 16'h1cb4, 16'h1cd0, 16'h1cec, 16'h1d08, 16'h1d24, 16'h1d40, 16'h1d5c, 16'h1d78, 16'h1d94, 16'h1db0, 16'h1dcc, 16'h1de8, 16'h1e04, 16'h1e20, 16'h1e3c, 16'h1e58, 16'h1e74, 16'h1e90, 16'h1eac, 16'h1ec8, 16'h1ee4, 16'h1f00, 16'h1f1c, 16'h1f38, 16'h1f54, 16'h1f70},
                                 {16'h1f8c, 16'h1fa8, 16'h1fc4, 16'h1fe0, 16'h1ffc, 16'h2018, 16'h2034, 16'h2050, 16'h206c, 16'h2088, 16'h20a4, 16'h20c0, 16'h20dc, 16'h20f8, 16'h2114, 16'h2130, 16'h214c, 16'h2168, 16'h2184, 16'h21a0, 16'h21bc, 16'h21d8, 16'h21f4, 16'h2210, 16'h222c, 16'h2248, 16'h2264, 16'h2280, 16'h229c, 16'h22b8, 16'h22d4, 16'h22f0, 16'h230c, 16'h2328, 16'h2344, 16'h2360, 16'h237c, 16'h2398, 16'h23b4, 16'h23d0, 16'h23ec, 16'h2408, 16'h2424, 16'h2440, 16'h245c, 16'h2478, 16'h2494, 16'h24b0, 16'h24cc, 16'h24e8, 16'h2504, 16'h2520, 16'h253c, 16'h2558, 16'h2574, 16'h2590, 16'h25ac, 16'h25c8, 16'h25e4, 16'h2600, 16'h261c, 16'h2638, 16'h2654, 16'h2670},
                                 {16'h268c, 16'h26a8, 16'h26c4, 16'h26e0, 16'h26fc, 16'h2718, 16'h2734, 16'h2750, 16'h276c, 16'h2788, 16'h27a4, 16'h27c0, 16'h27dc, 16'h27f8, 16'h2814, 16'h2830, 16'h284c, 16'h2868, 16'h2884, 16'h28a0, 16'h28bc, 16'h28d8, 16'h28f4, 16'h2910, 16'h292c, 16'h2948, 16'h2964, 16'h2980, 16'h299c, 16'h29b8, 16'h29d4, 16'h29f0, 16'h2a0c, 16'h2a28, 16'h2a44, 16'h2a60, 16'h2a7c, 16'h2a98, 16'h2ab4, 16'h2ad0, 16'h2aec, 16'h2b08, 16'h2b24, 16'h2b40, 16'h2b5c, 16'h2b78, 16'h2b94, 16'h2bb0, 16'h2bcc, 16'h2be8, 16'h2c04, 16'h2c20, 16'h2c3c, 16'h2c58, 16'h2c74, 16'h2c90, 16'h2cac, 16'h2cc8, 16'h2ce4, 16'h2d00, 16'h2d1c, 16'h2d38, 16'h2d54, 16'h2d70},
                                 {16'h2d8c, 16'h2da8, 16'h2dc4, 16'h2de0, 16'h2dfc, 16'h2e18, 16'h2e34, 16'h2e50, 16'h2e6c, 16'h2e88, 16'h2ea4, 16'h2ec0, 16'h2edc, 16'h2ef8, 16'h2f14, 16'h2f30, 16'h2f4c, 16'h2f68, 16'h2f84, 16'h2fa0, 16'h2fbc, 16'h2fd8, 16'h2ff4, 16'h3010, 16'h302c, 16'h3048, 16'h3064, 16'h3080, 16'h309c, 16'h30b8, 16'h30d4, 16'h30f0, 16'h310c, 16'h3128, 16'h3144, 16'h3160, 16'h317c, 16'h3198, 16'h31b4, 16'h31d0, 16'h31ec, 16'h3208, 16'h3224, 16'h3240, 16'h325c, 16'h3278, 16'h3294, 16'h32b0, 16'h32cc, 16'h32e8, 16'h3304, 16'h3320, 16'h333c, 16'h3358, 16'h3374, 16'h3390, 16'h33ac, 16'h33c8, 16'h33e4, 16'h3400, 16'h341c, 16'h3438, 16'h3454, 16'h3470},
                                 {16'h348c, 16'h34a8, 16'h34c4, 16'h34e0, 16'h34fc, 16'h3518, 16'h3534, 16'h3550, 16'h37bc, 16'h37bc, 16'h37bc, 16'h37bc, 16'h37bc, 16'h37bc, 16'h37bc, 16'h37bc, 16'h37bc, 16'h37bc, 16'h37bc, 16'h37bc, 16'h37bc, 16'h37bc, 16'h37bc, 16'h37bc, 16'h37bc, 16'h37bc, 16'h37bc, 16'h37bc, 16'h37bc, 16'h37b7, 16'h37b1, 16'h37ab, 16'h37a5, 16'h379f, 16'h3799, 16'h3793, 16'h378d, 16'h3787, 16'h3781, 16'h377b, 16'h3775, 16'h376f, 16'h3769, 16'h3763, 16'h375d, 16'h3757, 16'h3751, 16'h374b, 16'h3745, 16'h373f, 16'h3739, 16'h3733, 16'h372d, 16'h3727, 16'h3721, 16'h371b, 16'h3715, 16'h370f, 16'h3709, 16'h3703, 16'h36fd, 16'h36f7, 16'h36f1, 16'h36eb},
                                 {16'h36e5, 16'h36df, 16'h36d9, 16'h36d3, 16'h36cd, 16'h36c7, 16'h36c1, 16'h36bb, 16'h36b5, 16'h36af, 16'h36a9, 16'h36a3, 16'h369d, 16'h3697, 16'h3691, 16'h368b, 16'h3685, 16'h367f, 16'h3679, 16'h3673, 16'h366d, 16'h3667, 16'h3661, 16'h365b, 16'h3655, 16'h364f, 16'h3649, 16'h3643, 16'h363d, 16'h3637, 16'h3631, 16'h362b, 16'h3625, 16'h361f, 16'h3619, 16'h3613, 16'h360d, 16'h3607, 16'h3601, 16'h35fb, 16'h35f5, 16'h35ef, 16'h35e9, 16'h35e3, 16'h35dd, 16'h35d7, 16'h35d1, 16'h35cb, 16'h35c5, 16'h35bf, 16'h35b9, 16'h35b3, 16'h35ad, 16'h35a7, 16'h35a1, 16'h359b, 16'h3595, 16'h358f, 16'h3589, 16'h3583, 16'h357d, 16'h3577, 16'h3571, 16'h356b},
                                 {16'h3565, 16'h355f, 16'h3559, 16'h3553, 16'h354d, 16'h3547, 16'h3541, 16'h353b, 16'h3535, 16'h352f, 16'h3529, 16'h3523, 16'h351d, 16'h3517, 16'h3511, 16'h350b, 16'h3505, 16'h34ff, 16'h34f9, 16'h34f3, 16'h34ed, 16'h34e7, 16'h34e1, 16'h34db, 16'h34d5, 16'h34cf, 16'h34c9, 16'h34c3, 16'h34bd, 16'h34b7, 16'h34b1, 16'h34ab, 16'h34a5, 16'h349f, 16'h3499, 16'h3493, 16'h348d, 16'h3487, 16'h3481, 16'h347b, 16'h3475, 16'h346f, 16'h3469, 16'h3463, 16'h345d, 16'h3457, 16'h3451, 16'h344b, 16'h3445, 16'h343f, 16'h3439, 16'h3433, 16'h342d, 16'h3427, 16'h3421, 16'h341b, 16'h3415, 16'h340f, 16'h3409, 16'h3403, 16'h33fd, 16'h33f7, 16'h33f1, 16'h33eb},
                                 {16'h33e5, 16'h33df, 16'h33d9, 16'h33d3, 16'h33cd, 16'h33c7, 16'h33c1, 16'h33bb, 16'h33b5, 16'h33af, 16'h33a9, 16'h33a3, 16'h339d, 16'h3397, 16'h3391, 16'h338b, 16'h3385, 16'h337f, 16'h3379, 16'h3373, 16'h336d, 16'h3367, 16'h3361, 16'h335b, 16'h3355, 16'h334f, 16'h3349, 16'h3343, 16'h333d, 16'h3337, 16'h3331, 16'h332b, 16'h3325, 16'h331f, 16'h3319, 16'h3313, 16'h330d, 16'h3307, 16'h3301, 16'h32fb, 16'h32f5, 16'h32ef, 16'h32e9, 16'h32e3, 16'h32dd, 16'h32d7, 16'h32d1, 16'h32cb, 16'h32c5, 16'h32bf, 16'h32b9, 16'h32b3, 16'h32ad, 16'h32a7, 16'h32a1, 16'h329b, 16'h3295, 16'h328f, 16'h3289, 16'h3283, 16'h327d, 16'h3277, 16'h3271, 16'h326b},
                                 {16'h3265, 16'h325f, 16'h3259, 16'h3253, 16'h324d, 16'h3247, 16'h3241, 16'h323b, 16'h3235, 16'h322f, 16'h3229, 16'h3223, 16'h321d, 16'h3217, 16'h3211, 16'h320b, 16'h3205, 16'h31ff, 16'h31f9, 16'h31f3, 16'h31ed, 16'h31e7, 16'h31e1, 16'h31db, 16'h31d5, 16'h31cf, 16'h31c9, 16'h31c3, 16'h31bd, 16'h31b7, 16'h31b1, 16'h31ab, 16'h31a5, 16'h319f, 16'h3199, 16'h3193, 16'h318d, 16'h3187, 16'h3181, 16'h317b, 16'h3175, 16'h316f, 16'h3169, 16'h3163, 16'h315d, 16'h3157, 16'h3151, 16'h314b, 16'h3145, 16'h313f, 16'h3139, 16'h3133, 16'h312d, 16'h3127, 16'h3121, 16'h311b, 16'h3115, 16'h310f, 16'h3109, 16'h3103, 16'h30fd, 16'h30f7, 16'h30f1, 16'h30eb},
                                 {16'h30e5, 16'h30df, 16'h30d9, 16'h30d3, 16'h30cd, 16'h30c7, 16'h30c1, 16'h30bb, 16'h30b5, 16'h30af, 16'h30a9, 16'h30a3, 16'h309d, 16'h3097, 16'h3091, 16'h308b, 16'h3085, 16'h307f, 16'h3079, 16'h3073, 16'h306d, 16'h3067, 16'h3061, 16'h305b, 16'h3055, 16'h304f, 16'h3049, 16'h3043, 16'h303d, 16'h3037, 16'h3031, 16'h302b, 16'h3025, 16'h301f, 16'h3019, 16'h3013, 16'h300d, 16'h3007, 16'h3001, 16'h2ffb, 16'h2ff5, 16'h2fef, 16'h2fe9, 16'h2fe3, 16'h2fdd, 16'h2fd7, 16'h2fd1, 16'h2fcb, 16'h2fc5, 16'h2fbf, 16'h2fb9, 16'h2fb3, 16'h2fad, 16'h2fa7, 16'h2fa1, 16'h2f9b, 16'h2f95, 16'h2f8f, 16'h2f89, 16'h2f83, 16'h2f7d, 16'h2f77, 16'h2f71, 16'h2f6b},
                                 {16'h2f65, 16'h2f5f, 16'h2f59, 16'h2f53, 16'h2f4d, 16'h2f47, 16'h2f41, 16'h2f3b, 16'h2f35, 16'h2f2f, 16'h2f29, 16'h2f23, 16'h2f1d, 16'h2f17, 16'h2f11, 16'h2f0b, 16'h2f05, 16'h2eff, 16'h2ef9, 16'h2ef3, 16'h2eed, 16'h2ee7, 16'h2ee1, 16'h2edb, 16'h2ed5, 16'h2ecf, 16'h2ec9, 16'h2ec3, 16'h2ebd, 16'h2eb7, 16'h2eb1, 16'h2eab, 16'h2ea5, 16'h2e9f, 16'h2e99, 16'h2e93, 16'h2e8d, 16'h2e87, 16'h2e81, 16'h2e7b, 16'h2e75, 16'h2e6f, 16'h2e69, 16'h2e63, 16'h2e5d, 16'h2e57, 16'h2e51, 16'h2e4b, 16'h2e45, 16'h2e3f, 16'h2e39, 16'h2e33, 16'h2e2d, 16'h2e27, 16'h2e21, 16'h2e1b, 16'h2e15, 16'h2e0f, 16'h2e09, 16'h2e03, 16'h2dfd, 16'h2df7, 16'h2df1, 16'h2deb},
                                 {16'h2de5, 16'h2ddf, 16'h2dd9, 16'h2dd3, 16'h2dcd, 16'h2dc7, 16'h2dc1, 16'h2dbb, 16'h2db5, 16'h2daf, 16'h2da9, 16'h2da3, 16'h2d9d, 16'h2d97, 16'h2d91, 16'h2d8b, 16'h2d85, 16'h2d7f, 16'h2d79, 16'h2d73, 16'h2d6d, 16'h2d67, 16'h2d61, 16'h2d5b, 16'h2d55, 16'h2d4f, 16'h2d49, 16'h2d43, 16'h2d3d, 16'h2d37, 16'h2d31, 16'h2d2b, 16'h2d25, 16'h2d1f, 16'h2d19, 16'h2d13, 16'h2d0d, 16'h2d07, 16'h2d01, 16'h2cfb, 16'h2cf5, 16'h2cef, 16'h2ce9, 16'h2ce3, 16'h2cdd, 16'h2cd7, 16'h2cd1, 16'h2ccb, 16'h2cc5, 16'h2cbf, 16'h2cb9, 16'h2cb3, 16'h2cad, 16'h2ca7, 16'h2ca1, 16'h2c9b, 16'h2c95, 16'h2c8f, 16'h2c89, 16'h2c83, 16'h2c7d, 16'h2c77, 16'h2c71, 16'h2c6b},
                                 {16'h2c65, 16'h2c5f, 16'h2c59, 16'h2c53, 16'h2c4d, 16'h2c47, 16'h2c41, 16'h2c3b, 16'h2c35, 16'h2c2f, 16'h2c29, 16'h2c23, 16'h2c1d, 16'h2c17, 16'h2c11, 16'h2c0b, 16'h2c05, 16'h2bff, 16'h2bf9, 16'h2bf3, 16'h2bed, 16'h2be7, 16'h2be1, 16'h2bdb, 16'h2bd5, 16'h2bcf, 16'h2bc9, 16'h2bc3, 16'h2bbd, 16'h2bb7, 16'h2bb1, 16'h2bb1, 16'h2bb1, 16'h2bb1, 16'h2bb1, 16'h2baa, 16'h2b9b, 16'h2b8c, 16'h2b7d, 16'h2b6e, 16'h2b5f, 16'h2b50, 16'h2b41, 16'h2b32, 16'h2b23, 16'h2b14, 16'h2b05, 16'h2af6, 16'h2ae7, 16'h2ad8, 16'h2ac9, 16'h2aba, 16'h2aab, 16'h2a9c, 16'h2a8d, 16'h2a7e, 16'h2a6f, 16'h2a60, 16'h2a51, 16'h2a42, 16'h2a33, 16'h2a24, 16'h2a15, 16'h2a06},
                                 {16'h29f7, 16'h29e8, 16'h29d9, 16'h29ca, 16'h29bb, 16'h29ac, 16'h299d, 16'h298e, 16'h297f, 16'h2970, 16'h2961, 16'h2952, 16'h2943, 16'h2934, 16'h2925, 16'h2916, 16'h2907, 16'h28f8, 16'h28e9, 16'h28da, 16'h28cb, 16'h28bc, 16'h28ad, 16'h289e, 16'h288f, 16'h2880, 16'h2871, 16'h2862, 16'h2853, 16'h2844, 16'h2835, 16'h2826, 16'h2817, 16'h2808, 16'h27f9, 16'h27ea, 16'h27db, 16'h27cc, 16'h27bd, 16'h27ae, 16'h279f, 16'h2790, 16'h2781, 16'h2772, 16'h2763, 16'h2754, 16'h2745, 16'h2736, 16'h2727, 16'h2718, 16'h2709, 16'h26fa, 16'h26eb, 16'h26dc, 16'h26cd, 16'h26be, 16'h26af, 16'h26a0, 16'h2691, 16'h2682, 16'h2673, 16'h2664, 16'h2655, 16'h2646},
                                 {16'h2637, 16'h2628, 16'h2619, 16'h260a, 16'h25fb, 16'h25ec, 16'h25dd, 16'h25ce, 16'h25bf, 16'h25b0, 16'h25a1, 16'h2592, 16'h2583, 16'h2574, 16'h2565, 16'h2556, 16'h2547, 16'h2538, 16'h2529, 16'h251a, 16'h250b, 16'h24fc, 16'h24ed, 16'h24de, 16'h24cf, 16'h24c0, 16'h24b1, 16'h24a2, 16'h2493, 16'h2484, 16'h2475, 16'h2466, 16'h2457, 16'h2448, 16'h2439, 16'h242a, 16'h241b, 16'h240c, 16'h23fd, 16'h23ee, 16'h23df, 16'h23d0, 16'h23c1, 16'h23b2, 16'h23a3, 16'h2394, 16'h2385, 16'h2376, 16'h2367, 16'h2358, 16'h2349, 16'h233a, 16'h232b, 16'h231c, 16'h230d, 16'h22fe, 16'h22ef, 16'h22e0, 16'h2316, 16'h234a, 16'h237e, 16'h23b2, 16'h23e6, 16'h241a},
                                 {16'h244e, 16'h2482, 16'h24b6, 16'h24ea, 16'h251e, 16'h2552, 16'h2586, 16'h25ba, 16'h25ee, 16'h2622, 16'h2557, 16'h253f, 16'h2527, 16'h250f, 16'h24f7, 16'h24df, 16'h24c7, 16'h24af, 16'h2497, 16'h247f, 16'h2467, 16'h244f, 16'h2437, 16'h241f, 16'h2407, 16'h23ef, 16'h23d7, 16'h23bf, 16'h23a7, 16'h238f, 16'h2377, 16'h235f, 16'h2347, 16'h232f, 16'h2317, 16'h22ff, 16'h22e7, 16'h22cf, 16'h22b7, 16'h229f, 16'h2287, 16'h226f, 16'h2257, 16'h223f, 16'h2227, 16'h220f, 16'h21f7, 16'h21df, 16'h21c7, 16'h21af, 16'h2197, 16'h217f, 16'h2167, 16'h214f, 16'h2137, 16'h211f, 16'h2107, 16'h20ef, 16'h20d7, 16'h20bf, 16'h20a7, 16'h208f, 16'h2077, 16'h205f},
                                 {16'h2047, 16'h202f, 16'h2017, 16'h1fff, 16'h1fe7, 16'h1fcf, 16'h1fb7, 16'h1f9f, 16'h1f87, 16'h1f6f, 16'h1f57, 16'h1f3f, 16'h1f27, 16'h1f0f, 16'h1ef7, 16'h1edf, 16'h1ec7, 16'h1eaf, 16'h1e97, 16'h1e7f, 16'h1e67, 16'h1e4f, 16'h1e37, 16'h1e1f, 16'h1e07, 16'h1def, 16'h1dd7, 16'h1dbf, 16'h1da7, 16'h1d8f, 16'h1d77, 16'h1d5f, 16'h1d47, 16'h1d2f, 16'h1d17, 16'h1cff, 16'h1ce7, 16'h1ccf, 16'h1cb7, 16'h1c9f, 16'h1c87, 16'h1c6f, 16'h1c57, 16'h1c3f, 16'h1c27, 16'h1c0f, 16'h1bf7, 16'h1bdf, 16'h1bc7, 16'h1baf, 16'h1b97, 16'h1b7f, 16'h1b67, 16'h1b4f, 16'h1b37, 16'h1b1f, 16'h1b07, 16'h1aef, 16'h1ad7, 16'h1abf, 16'h1aa7, 16'h1a8f, 16'h1a77, 16'h1a5f},
                                 {16'h1a47, 16'h1a2f, 16'h1a17, 16'h19ff, 16'h19e7, 16'h19cf, 16'h19b7, 16'h199f, 16'h1987, 16'h196f, 16'h1957, 16'h193f, 16'h1927, 16'h190f, 16'h18f7, 16'h18df, 16'h18c7, 16'h18af, 16'h1897, 16'h187f, 16'h1867, 16'h184f, 16'h1837, 16'h181f, 16'h1807, 16'h17ef, 16'h17d7, 16'h17bf, 16'h17a7, 16'h178f, 16'h1777, 16'h175f, 16'h1747, 16'h172f, 16'h1717, 16'h16ff, 16'h16e7, 16'h16cf, 16'h16b7, 16'h169f, 16'h1687, 16'h166f, 16'h1657, 16'h163f, 16'h1627, 16'h160f, 16'h15f7, 16'h15df, 16'h15c7, 16'h15af, 16'h1597, 16'h157f, 16'h1567, 16'h154f, 16'h1537, 16'h151f, 16'h1507, 16'h14ef, 16'h14d7, 16'h14bf, 16'h14a7, 16'h148f, 16'h1477, 16'h145f},
                                 {16'h1447, 16'h142f, 16'h1417, 16'h13ff, 16'h13e7, 16'h13cf, 16'h13b7, 16'h139f, 16'h1387, 16'h136f, 16'h1357, 16'h133f, 16'h1327, 16'h130f, 16'h12f7, 16'h12df, 16'h12c7, 16'h12af, 16'h1297, 16'h127f, 16'h1267, 16'h124f, 16'h1237, 16'h121f, 16'h1207, 16'h11ef, 16'h11d7, 16'h11bf, 16'h11a7, 16'h118f, 16'h1177, 16'h115f, 16'h1147, 16'h112f, 16'h1117, 16'h10ff, 16'h10e7, 16'h10cf, 16'h10b7, 16'h109f, 16'h1087, 16'h106f, 16'h1057, 16'h103f, 16'h1027, 16'h100f, 16'h0ff7, 16'h0fdf, 16'h0fc7, 16'h0faf, 16'h0f97, 16'h0f7f, 16'h0f67, 16'h0f4f, 16'h0f37, 16'h0f1f, 16'h0f07, 16'h0eef, 16'h0ed7, 16'h0ebf, 16'h0ea7, 16'h0e8f, 16'h0e77, 16'h0e5f},
                                 {16'h0e47, 16'h0e2f, 16'h0e17, 16'h0dff, 16'h0de7, 16'h0dcf, 16'h0db7, 16'h0d9f, 16'h0d87, 16'h0d6f, 16'h0d57, 16'h0d3f, 16'h0d27, 16'h0d0f, 16'h0cf7, 16'h0cdf, 16'h0cc7, 16'h0caf, 16'h0c97, 16'h0c7f, 16'h0c67, 16'h0c4f, 16'h0c37, 16'h0c1f, 16'h0c07, 16'h0bef, 16'h0bd7, 16'h0bbf, 16'h0ba7, 16'h0b8f, 16'h0b77, 16'h0b5f, 16'h0b47, 16'h0b2f, 16'h0b17, 16'h0aff, 16'h0ae7, 16'h0acf, 16'h0ab7, 16'h0a9f, 16'h0a87, 16'h0a6f, 16'h0a57, 16'h0a3f, 16'h0a27, 16'h0a0f, 16'h09f7, 16'h09df, 16'h09c7, 16'h09af, 16'h0997, 16'h097f, 16'h0967, 16'h094f, 16'h0937, 16'h091f, 16'h0907, 16'h08ef, 16'h08d7, 16'h08bf, 16'h08a7, 16'h088f, 16'h0877, 16'h085f},
                                 {16'h0847, 16'h082f, 16'h0817, 16'h07ff, 16'h07e7, 16'h07cf, 16'h07b7, 16'h079f, 16'h0787, 16'h076f, 16'h0757, 16'h073f, 16'h0727, 16'h070f, 16'h06f7, 16'h06df, 16'h06c7, 16'h06af, 16'h0697, 16'h067f, 16'h0667, 16'h064f, 16'h0637, 16'h061f, 16'h0607, 16'h05ef, 16'h05d7, 16'h05bf, 16'h05a7, 16'h058f, 16'h0577, 16'h055f, 16'h0547, 16'h052f, 16'h0517, 16'h04ff, 16'h04e7, 16'h04cf, 16'h04b7, 16'h049f, 16'h0487, 16'h046f, 16'h0457, 16'h043f, 16'h0427, 16'h040f, 16'h03f7, 16'h03df, 16'h03c7, 16'h03af, 16'h0397, 16'h037f, 16'h0367, 16'h034f, 16'h0337, 16'h031f, 16'h0307, 16'h02ef, 16'h02d7, 16'h02bf, 16'h02a7, 16'h0349, 16'h03fa, 16'h04ab},
                                 {16'h055c, 16'h060d, 16'h06be, 16'h076f, 16'h0820, 16'h08d1, 16'h0982, 16'h0a33, 16'h0ae4, 16'h0b95, 16'h0c46, 16'h0cf7, 16'h0da8, 16'h0e59, 16'h0f0a, 16'h0fbb, 16'h106c, 16'h111d, 16'h11ce, 16'h127f, 16'h1330, 16'h13e1, 16'h1492, 16'h1543, 16'h15f4, 16'h16a5, 16'h1756, 16'h1807, 16'h18b8, 16'h1969, 16'h1a1a, 16'h1acb, 16'h1b7c, 16'h1c2d, 16'h1cde, 16'h1d8f, 16'h1e40, 16'h1ef1, 16'h1fa2, 16'h2053, 16'h2104, 16'h21b5, 16'h2266, 16'h2317, 16'h23c8, 16'h2479, 16'h2479, 16'h2479, 16'h2479, 16'h2479, 16'h2479, 16'h2479, 16'h2479, 16'h246d, 16'h245d, 16'h244d, 16'h243d, 16'h242d, 16'h241d, 16'h240d, 16'h23fd, 16'h23ed, 16'h23dd, 16'h23cd},
                                 {16'h23bd, 16'h23ad, 16'h239d, 16'h238d, 16'h237d, 16'h236d, 16'h235d, 16'h234d, 16'h233d, 16'h232d, 16'h231d, 16'h230d, 16'h22fd, 16'h22ed, 16'h22dd, 16'h22cd, 16'h22bd, 16'h22ad, 16'h229d, 16'h228d, 16'h227d, 16'h226d, 16'h225d, 16'h224d, 16'h223d, 16'h222d, 16'h221d, 16'h220d, 16'h21fd, 16'h21ed, 16'h21dd, 16'h21cd, 16'h21bd, 16'h21ad, 16'h219d, 16'h218d, 16'h217d, 16'h216d, 16'h215d, 16'h214d, 16'h213d, 16'h212d, 16'h211d, 16'h210d, 16'h20fd, 16'h20ed, 16'h20dd, 16'h20cd, 16'h20bd, 16'h20ad, 16'h209d, 16'h208d, 16'h207d, 16'h206d, 16'h205d, 16'h204d, 16'h203d, 16'h202d, 16'h201d, 16'h200d, 16'h1ffd, 16'h1fed, 16'h1fdd, 16'h1fcd},
                                 {16'h1fbd, 16'h1fad, 16'h1f9d, 16'h1f8d, 16'h1f7d, 16'h1f6d, 16'h1f5d, 16'h1f4d, 16'h1f3d, 16'h1f2d, 16'h1f1d, 16'h1f0d, 16'h1efd, 16'h1eed, 16'h1edd, 16'h1ecd, 16'h1ebd, 16'h1ead, 16'h1e9d, 16'h1e8d, 16'h1e7d, 16'h1e6d, 16'h1e5d, 16'h1e4d, 16'h1e3d, 16'h1e2d, 16'h1e1d, 16'h1e0d, 16'h1dfd, 16'h1ded, 16'h1ddd, 16'h1dcd, 16'h1dbd, 16'h1dad, 16'h1d9d, 16'h1d8d, 16'h1d7d, 16'h1d6d, 16'h1d5d, 16'h1d4d, 16'h1d3d, 16'h1d2d, 16'h1d1d, 16'h1d0d, 16'h1cfd, 16'h1ced, 16'h1cdd, 16'h1ccd, 16'h1cbd, 16'h1cad, 16'h1c9d, 16'h1c8d, 16'h1c7d, 16'h1c6d, 16'h1c5d, 16'h1c4d, 16'h1c3d, 16'h1c2d, 16'h1c1d, 16'h1c0d, 16'h1bfd, 16'h1bed, 16'h1bdd, 16'h1bcd},
                                 {16'h1bbd, 16'h1bad, 16'h1b9d, 16'h1b8d, 16'h1b7d, 16'h1b6d, 16'h1b5d, 16'h1b4d, 16'h1b3d, 16'h1b2d, 16'h1b1d, 16'h1b0d, 16'h1afd, 16'h1aed, 16'h1add, 16'h1acd, 16'h1abd, 16'h1aad, 16'h1a9d, 16'h1a8d, 16'h1a7d, 16'h1a6d, 16'h1a5d, 16'h1a4d, 16'h1a3d, 16'h1a2d, 16'h1a1d, 16'h1a0d, 16'h19fd, 16'h19ed, 16'h19dd, 16'h19cd, 16'h19bd, 16'h19ad, 16'h199d, 16'h198d, 16'h197d, 16'h196d, 16'h195d, 16'h194d, 16'h193d, 16'h192d, 16'h191d, 16'h190d, 16'h18fd, 16'h18ed, 16'h18dd, 16'h18cd, 16'h18bd, 16'h18ad, 16'h189d, 16'h188d, 16'h187d, 16'h186d, 16'h185d, 16'h184d, 16'h183d, 16'h182d, 16'h181d, 16'h180d, 16'h17fd, 16'h17ed, 16'h17dd, 16'h17cd},
                                 {16'h17bd, 16'h17ad, 16'h179d, 16'h178d, 16'h177d, 16'h176d, 16'h175d, 16'h174d, 16'h173d, 16'h172d, 16'h171d, 16'h170d, 16'h16fd, 16'h16ed, 16'h16dd, 16'h16cd, 16'h16bd, 16'h16ad, 16'h169d, 16'h168d, 16'h167d, 16'h166d, 16'h165d, 16'h164d, 16'h163d, 16'h162d, 16'h161d, 16'h160d, 16'h15fd, 16'h15ed, 16'h15dd, 16'h15cd, 16'h15bd, 16'h15ad, 16'h159d, 16'h158d, 16'h157d, 16'h156d, 16'h155d, 16'h154d, 16'h153d, 16'h152d, 16'h151d, 16'h150d, 16'h14fd, 16'h14ed, 16'h14dd, 16'h14cd, 16'h14bd, 16'h14ad, 16'h149d, 16'h148d, 16'h147d, 16'h146d, 16'h145d, 16'h144d, 16'h143d, 16'h142d, 16'h141d, 16'h140d, 16'h13fd, 16'h13ed, 16'h13dd, 16'h13cd},
                                 {16'h13bd, 16'h13ad, 16'h139d, 16'h138d, 16'h137d, 16'h136d, 16'h135d, 16'h134d, 16'h133d, 16'h132d, 16'h131d, 16'h130d, 16'h12fd, 16'h12ed, 16'h12dd, 16'h12cd, 16'h12bd, 16'h12ad, 16'h129d, 16'h128d, 16'h127d, 16'h126d, 16'h125d, 16'h124d, 16'h123d, 16'h122d, 16'h121d, 16'h120d, 16'h11fd, 16'h11ed, 16'h11dd, 16'h11cd, 16'h11bd, 16'h11ad, 16'h119d, 16'h118d, 16'h117d, 16'h116d, 16'h115d, 16'h114d, 16'h113d, 16'h112d, 16'h111d, 16'h110d, 16'h10fd, 16'h10ed, 16'h10dd, 16'h10cd, 16'h10bd, 16'h10ad, 16'h109d, 16'h108d, 16'h107d, 16'h106d, 16'h105d, 16'h104d, 16'h103d, 16'h102d, 16'h101d, 16'h100d, 16'h0ffd, 16'h0fed, 16'h0fdd, 16'h0fcd},
                                 {16'h0fbd, 16'h0fad, 16'h0f9d, 16'h0f8d, 16'h0f7d, 16'h0f6d, 16'h0f5d, 16'h0f4d, 16'h0f3d, 16'h0f2d, 16'h0f1d, 16'h0f0d, 16'h0efd, 16'h0eed, 16'h0edd, 16'h0ecd, 16'h0ebd, 16'h0ead, 16'h0e9d, 16'h0e8d, 16'h0e7d, 16'h0e6d, 16'h0e5d, 16'h0e4d, 16'h0e3d, 16'h0e2d, 16'h0e1d, 16'h0e0d, 16'h0dfd, 16'h0ded, 16'h0ddd, 16'h0dcd, 16'h0dbd, 16'h0dad, 16'h0d9d, 16'h0d8d, 16'h0d7d, 16'h0d6d, 16'h0d5d, 16'h0d4d, 16'h0d3d, 16'h0d2d, 16'h0d1d, 16'h0d0d, 16'h0cfd, 16'h0ced, 16'h0cdd, 16'h0ccd, 16'h0cbd, 16'h0cad, 16'h0c9d, 16'h0c8d, 16'h0c7d, 16'h0c6d, 16'h0c5d, 16'h0c4d, 16'h0c3d, 16'h0c2d, 16'h0c1d, 16'h0c0d, 16'h0bfd, 16'h0bed, 16'h0bdd, 16'h0bcd},
                                 {16'h0bbd, 16'h0bad, 16'h0b9d, 16'h0b8d, 16'h0b7d, 16'h0b6d, 16'h0b62, 16'h0b61, 16'h0b60, 16'h0b5f, 16'h0b5e, 16'h0b5d, 16'h0b5c, 16'h0b5b, 16'h0b5a, 16'h0b59, 16'h0b58, 16'h0b57, 16'h0b56, 16'h0b55, 16'h0b54, 16'h0b53, 16'h0b52, 16'h0b51, 16'h0b50, 16'h0b4f, 16'h0b4e, 16'h0b4d, 16'h0b4c, 16'h0b4b, 16'h0b4a, 16'h0b49, 16'h0b48, 16'h0b47, 16'h0b46, 16'h0b45, 16'h0b44, 16'h0b43, 16'h0b42, 16'h0b41, 16'h0b40, 16'h0b3f, 16'h0b3e, 16'h0b3d, 16'h0b3c, 16'h0b3b, 16'h0b3a, 16'h0b39, 16'h0b38, 16'h0b37, 16'h0b36, 16'h0b35, 16'h0b34, 16'h0b33, 16'h0b32, 16'h0b31, 16'h0b30, 16'h0b2f, 16'h0b2e, 16'h0b2d, 16'h0b2c, 16'h0b2b, 16'h0b2a, 16'h0b29},
                                 {16'h0b28, 16'h0b27, 16'h0b26, 16'h0b25, 16'h0b24, 16'h0b23, 16'h0b22, 16'h0b21, 16'h0b20, 16'h0b1f, 16'h0b1e, 16'h0b1d, 16'h0b1c, 16'h0b1b, 16'h0b1a, 16'h0b19, 16'h0b18, 16'h0b17, 16'h0b16, 16'h0b15, 16'h0b14, 16'h0b13, 16'h0b12, 16'h0b11, 16'h0b10, 16'h0b0f, 16'h0b0e, 16'h0b0d, 16'h0b0c, 16'h0b0b, 16'h0b0a, 16'h0b09, 16'h0b08, 16'h0b07, 16'h0b06, 16'h0b05, 16'h0b04, 16'h0b03, 16'h0b02, 16'h0b01, 16'h0b00, 16'h0aff, 16'h0afe, 16'h0afd, 16'h0afc, 16'h0afb, 16'h0afa, 16'h0af9, 16'h0af8, 16'h0af7, 16'h0af6, 16'h0af5, 16'h0af4, 16'h0af3, 16'h0af2, 16'h0af1, 16'h0af0, 16'h0aef, 16'h0aee, 16'h0aed, 16'h0aec, 16'h0aeb, 16'h0aea, 16'h0ae9},
                                 {16'h0ae8, 16'h0ae7, 16'h0ae6, 16'h0ae5, 16'h0ae4, 16'h0ae3, 16'h0ae2, 16'h0ae1, 16'h0ae0, 16'h0adf, 16'h0ade, 16'h0add, 16'h0adc, 16'h0adb, 16'h0ada, 16'h0ad9, 16'h0ad8, 16'h0ad7, 16'h0ad6, 16'h0ad5, 16'h0ad4, 16'h0ad3, 16'h0ad2, 16'h0ad1, 16'h0ad0, 16'h0acf, 16'h0ace, 16'h0acd, 16'h0acc, 16'h0acb, 16'h0aca, 16'h0ac9, 16'h0ac8, 16'h0ac7, 16'h0ac6, 16'h0ac5, 16'h0ac4, 16'h0ac3, 16'h0ac2, 16'h0ac1, 16'h0ac0, 16'h0abf, 16'h0abe, 16'h0abd, 16'h0abc, 16'h0abb, 16'h0aba, 16'h0ab9, 16'h0ab8, 16'h0ab7, 16'h0ab6, 16'h0ab5, 16'h0ab4, 16'h0ab3, 16'h0ab2, 16'h0ab1, 16'h0ab0, 16'h0aaf, 16'h0aae, 16'h0aad, 16'h0aac, 16'h0aab, 16'h0aaa, 16'h0aa9},
                                 {16'h0aa8, 16'h0aa7, 16'h0aa6, 16'h0aa5, 16'h0aa4, 16'h0aa3, 16'h0aa2, 16'h0aa1, 16'h0aa0, 16'h0a9f, 16'h0a9e, 16'h0a9d, 16'h0a9c, 16'h0a9b, 16'h0a9a, 16'h0a99, 16'h0a98, 16'h0a97, 16'h0a96, 16'h0a95, 16'h0a94, 16'h0a93, 16'h0a92, 16'h0a91, 16'h0a90, 16'h0b04, 16'h0b20, 16'h0b3c, 16'h0b58, 16'h0b74, 16'h0b90, 16'h0bac, 16'h0bc8, 16'h0be4, 16'h0c00, 16'h0c1c, 16'h0c38, 16'h0c54, 16'h0c70, 16'h0c8c, 16'h0ca8, 16'h0cc4, 16'h0ce0, 16'h0cfc, 16'h0d18, 16'h0d34, 16'h0d50, 16'h0d6c, 16'h0d88, 16'h0da4, 16'h0dc0, 16'h0ddc, 16'h0df8, 16'h0e14, 16'h0e30, 16'h0e4c, 16'h0e68, 16'h0e84, 16'h0ea0, 16'h0ebc, 16'h0ed8, 16'h0ef4, 16'h0f10, 16'h0f2c},
                                 {16'h0f48, 16'h0f64, 16'h0f80, 16'h0f9c, 16'h0fb8, 16'h0fd4, 16'h0ff0, 16'h100c, 16'h1028, 16'h1044, 16'h1060, 16'h107c, 16'h1098, 16'h10b4, 16'h10d0, 16'h10ec, 16'h1108, 16'h1124, 16'h1140, 16'h115c, 16'h1178, 16'h1194, 16'h11b0, 16'h11cc, 16'h11e8, 16'h1204, 16'h1220, 16'h123c, 16'h1258, 16'h1274, 16'h1290, 16'h12ac, 16'h12c8, 16'h12e4, 16'h1300, 16'h131c, 16'h1338, 16'h1354, 16'h1370, 16'h138c, 16'h13a8, 16'h13c4, 16'h13e0, 16'h13fc, 16'h1418, 16'h1434, 16'h1450, 16'h146c, 16'h1488, 16'h14a4, 16'h14c0, 16'h14dc, 16'h14f8, 16'h1514, 16'h1530, 16'h154c, 16'h1568, 16'h1584, 16'h15a0, 16'h15bc, 16'h15d8, 16'h15f4, 16'h1610, 16'h162c},
                                 {16'h1648, 16'h1664, 16'h1680, 16'h169c, 16'h16b8, 16'h16d4, 16'h16f0, 16'h170c, 16'h1728, 16'h1744, 16'h1760, 16'h177c, 16'h1798, 16'h17b4, 16'h17d0, 16'h17ec, 16'h1808, 16'h1824, 16'h1840, 16'h185c, 16'h1878, 16'h1894, 16'h18b0, 16'h18cc, 16'h18e8, 16'h1904, 16'h1920, 16'h193c, 16'h1958, 16'h1974, 16'h1990, 16'h19ac, 16'h19c8, 16'h19e4, 16'h1a00, 16'h1a1c, 16'h1a38, 16'h1a54, 16'h1a70, 16'h1a8c, 16'h1aa8, 16'h1ac4, 16'h1ae0, 16'h1afc, 16'h1b18, 16'h1b34, 16'h1b50, 16'h1b6c, 16'h1b88, 16'h1ba4, 16'h1bc0, 16'h1bdc, 16'h1bf8, 16'h1c14, 16'h1c30, 16'h1c4c, 16'h1c68, 16'h1c84, 16'h1ca0, 16'h1cbc, 16'h1cd8, 16'h1cf4, 16'h1d10, 16'h1d2c},
                                 {16'h1d48, 16'h1d64, 16'h1d80, 16'h1d9c, 16'h1db8, 16'h1dd4, 16'h1df0, 16'h1e0c, 16'h1e28, 16'h1e44, 16'h1e60, 16'h1e7c, 16'h1e98, 16'h1eb4, 16'h1ed0, 16'h1eec, 16'h1f08, 16'h1f24, 16'h1f40, 16'h1f5c, 16'h1f78, 16'h1f94, 16'h1fb0, 16'h1fcc, 16'h1fe8, 16'h2004, 16'h2020, 16'h203c, 16'h2058, 16'h2074, 16'h2090, 16'h20ac, 16'h20c8, 16'h20e4, 16'h2100, 16'h211c, 16'h2138, 16'h2154, 16'h2170, 16'h218c, 16'h21a8, 16'h21c4, 16'h21e0, 16'h21fc, 16'h2218, 16'h2234, 16'h2250, 16'h226c, 16'h2288, 16'h22a4, 16'h22c0, 16'h22dc, 16'h22f8, 16'h2314, 16'h2330, 16'h234c, 16'h2368, 16'h2384, 16'h23a0, 16'h23bc, 16'h23d8, 16'h23f4, 16'h2410, 16'h242c},
                                 {16'h2448, 16'h2464, 16'h2480, 16'h249c, 16'h24b8, 16'h24d4, 16'h24f0, 16'h250c, 16'h2528, 16'h2544, 16'h2560, 16'h257c, 16'h2598, 16'h25b4, 16'h25d0, 16'h25ec, 16'h2608, 16'h2624, 16'h2640, 16'h265c, 16'h2678, 16'h2694, 16'h26b0, 16'h26cc, 16'h26e8, 16'h2704, 16'h2720, 16'h273c, 16'h2758, 16'h2774, 16'h2790, 16'h27ac, 16'h27c8, 16'h27e4, 16'h2800, 16'h281c, 16'h2838, 16'h2854, 16'h2870, 16'h288c, 16'h28a8, 16'h28c4, 16'h28e0, 16'h28fc, 16'h2918, 16'h2934, 16'h2950, 16'h296c, 16'h2988, 16'h29a4, 16'h29c0, 16'h29dc, 16'h29f8, 16'h07bb, 16'h07bb, 16'h07bb, 16'h07bb, 16'h07db, 16'h0802, 16'h0829, 16'h0850, 16'h0877, 16'h089e, 16'h08c5},
                                 {16'h08ec, 16'h0913, 16'h093a, 16'h0961, 16'h0988, 16'h09af, 16'h09d6, 16'h09fd, 16'h0a24, 16'h0a4b, 16'h0a72, 16'h0a99, 16'h0ac0, 16'h0ae7, 16'h0b0e, 16'h0b35, 16'h0b5c, 16'h0b83, 16'h0baa, 16'h0bd1, 16'h0bf8, 16'h0c1f, 16'h0c46, 16'h0c6d, 16'h0c94, 16'h0cbb, 16'h0ce2, 16'h0d09, 16'h0d30, 16'h0d57, 16'h0d7e, 16'h0da5, 16'h0dcc, 16'h0df3, 16'h0e1a, 16'h0e41, 16'h0e68, 16'h0e8f, 16'h0eb6, 16'h0edd, 16'h0f04, 16'h0f2b, 16'h0f52, 16'h0f79, 16'h0fa0, 16'h0fc7, 16'h0fee, 16'h1015, 16'h103c, 16'h1063, 16'h108a, 16'h10b1, 16'h10d8, 16'h10ff, 16'h1126, 16'h114d, 16'h1174, 16'h119b, 16'h11c2, 16'h11e9, 16'h1210, 16'h1237, 16'h125e, 16'h1285},
                                 {16'h12ac, 16'h12d3, 16'h12fa, 16'h1321, 16'h1348, 16'h136f, 16'h1396, 16'h13bd, 16'h13e4, 16'h140b, 16'h1432, 16'h1459, 16'h1480, 16'h14a7, 16'h14ce, 16'h14f5, 16'h151c, 16'h1543, 16'h156a, 16'h1591, 16'h15b8, 16'h15df, 16'h1606, 16'h162d, 16'h1654, 16'h167b, 16'h16a2, 16'h16c9, 16'h16f0, 16'h1717, 16'h173e, 16'h1765, 16'h178c, 16'h17b3, 16'h17da, 16'h1801, 16'h1828, 16'h184f, 16'h1876, 16'h189d, 16'h18c4, 16'h18eb, 16'h1912, 16'h1939, 16'h1960, 16'h1987, 16'h19ae, 16'h19d5, 16'h19fc, 16'h1a23, 16'h1a4a, 16'h1a71, 16'h1a98, 16'h1abf, 16'h1ae6, 16'h1b0d, 16'h1b34, 16'h1b5b, 16'h1b82, 16'h1ba9, 16'h1bd0, 16'h1bf7, 16'h1c1e, 16'h1c45},
                                 {16'h1c6c, 16'h1c93, 16'h1cba, 16'h1ce1, 16'h1d08, 16'h1d2f, 16'h1d56, 16'h1d7d, 16'h1da4, 16'h1dcb, 16'h1df2, 16'h1e19, 16'h1e40, 16'h1e67, 16'h1e8e, 16'h1eb5, 16'h1edc, 16'h1f03, 16'h1f2a, 16'h1f51, 16'h1f78, 16'h1f9f, 16'h1fc6, 16'h1fed, 16'h2014, 16'h203b, 16'h2062, 16'h2089, 16'h20b0, 16'h20d7, 16'h20fe, 16'h2125, 16'h214c, 16'h2173, 16'h219a, 16'h21c1, 16'h21e8, 16'h220f, 16'h2236, 16'h225d, 16'h2284, 16'h22ab, 16'h22d2, 16'h22f9, 16'h2320, 16'h2347, 16'h236e, 16'h2395, 16'h23bc, 16'h23e3, 16'h240a, 16'h2431, 16'h2458, 16'h247f, 16'h24a6, 16'h24cd, 16'h24f4, 16'h251b, 16'h2542, 16'h2569, 16'h2590, 16'h25b7, 16'h25de, 16'h2605},
                                 {16'h262c, 16'h2653, 16'h267a, 16'h26a1, 16'h26c8, 16'h26ef, 16'h2716, 16'h273d, 16'h2764, 16'h278b, 16'h27b2, 16'h27d9, 16'h2800, 16'h2827, 16'h284e, 16'h2875, 16'h289c, 16'h28c3, 16'h28ea, 16'h2911, 16'h2938, 16'h295f, 16'h2986, 16'h29ad, 16'h29d4, 16'h29fb, 16'h2a22, 16'h2a49, 16'h2a70, 16'h2a97, 16'h2abe, 16'h2ae5, 16'h2b0c, 16'h2b33, 16'h2b5a, 16'h2b81, 16'h2ba8, 16'h2bcf, 16'h2bf6, 16'h2c1d, 16'h2c44, 16'h2c6b, 16'h2c92, 16'h2cb9, 16'h2ce0, 16'h2d07, 16'h2d2e, 16'h2d55, 16'h2d7c, 16'h2da3, 16'h2dca, 16'h2df1, 16'h2e18, 16'h2e3f, 16'h2e66, 16'h2e8d, 16'h2eb4, 16'h2edb, 16'h2f02, 16'h2f29, 16'h2f50, 16'h2f77, 16'h2f9e, 16'h2fc5},
                                 {16'h2fec, 16'h3013, 16'h303a, 16'h3061, 16'h3088, 16'h30af, 16'h30d6, 16'h30fd, 16'h3124, 16'h314b, 16'h3172, 16'h3199, 16'h31c0, 16'h31e7, 16'h320e, 16'h3235, 16'h325c, 16'h3283, 16'h32aa, 16'h32d1, 16'h32f8, 16'h331f, 16'h3346, 16'h336d, 16'h3394, 16'h33bb, 16'h33e2, 16'h3409, 16'h3430, 16'h3457, 16'h347e, 16'h34a5, 16'h34cc, 16'h34f3, 16'h351a, 16'h3541, 16'h3568, 16'h358f, 16'h35b6, 16'h35dd, 16'h3604, 16'h362b, 16'h3652, 16'h3679, 16'h36a0, 16'h36c7, 16'h36ee, 16'h3715, 16'h373c, 16'h3763, 16'h378a, 16'h37b1, 16'h37d8, 16'h37ff, 16'h3826, 16'h384d, 16'h3874, 16'h389b, 16'h38c2, 16'h38e9, 16'h3910, 16'h3937, 16'h3937, 16'h3937},
                                 {16'h3937, 16'h3925, 16'h3912, 16'h38ff, 16'h38ec, 16'h38d9, 16'h38c6, 16'h38b3, 16'h38a0, 16'h388d, 16'h387a, 16'h3867, 16'h3854, 16'h3841, 16'h382e, 16'h381b, 16'h3808, 16'h37f5, 16'h37e2, 16'h37cf, 16'h37bc, 16'h37a9, 16'h3796, 16'h3783, 16'h3770, 16'h375d, 16'h374a, 16'h3737, 16'h3724, 16'h3711, 16'h36fe, 16'h36eb, 16'h36d8, 16'h36c5, 16'h36b2, 16'h369f, 16'h368c, 16'h3679, 16'h3666, 16'h3653, 16'h3640, 16'h362d, 16'h361a, 16'h3607, 16'h35f4, 16'h35e1, 16'h35ce, 16'h35bb, 16'h35a8, 16'h3595, 16'h3582, 16'h356f, 16'h355c, 16'h3549, 16'h3536, 16'h3523, 16'h3510, 16'h34fd, 16'h34ea, 16'h34d7, 16'h34c4, 16'h34b1, 16'h349e, 16'h348b},
                                 {16'h3478, 16'h3465, 16'h3452, 16'h343f, 16'h342c, 16'h3419, 16'h3406, 16'h33f3, 16'h33e0, 16'h33cd, 16'h33ba, 16'h33a7, 16'h3394, 16'h3381, 16'h336e, 16'h335b, 16'h3348, 16'h3335, 16'h3322, 16'h330f, 16'h32fc, 16'h32e9, 16'h32d6, 16'h32c3, 16'h32b0, 16'h329d, 16'h328a, 16'h3277, 16'h3264, 16'h3251, 16'h323e, 16'h322b, 16'h3218, 16'h3205, 16'h31f2, 16'h31df, 16'h31cc, 16'h31b9, 16'h31a6, 16'h3193, 16'h3180, 16'h316d, 16'h315a, 16'h3147, 16'h3134, 16'h3121, 16'h310e, 16'h30fb, 16'h30e8, 16'h30d5, 16'h30c2, 16'h30af, 16'h309c, 16'h3089, 16'h3076, 16'h3063, 16'h3050, 16'h303d, 16'h302a, 16'h3017, 16'h3004, 16'h2ff1, 16'h2fde, 16'h2fcb},
                                 {16'h2fb8, 16'h2fa5, 16'h2f92, 16'h2f7f, 16'h2f6c, 16'h2f59, 16'h2f46, 16'h2f33, 16'h2f20, 16'h2f0d, 16'h2efa, 16'h2ee7, 16'h2ed4, 16'h2ec1, 16'h2eae, 16'h2e9b, 16'h2e88, 16'h2e75, 16'h2e62, 16'h2e4f, 16'h2e3c, 16'h2e29, 16'h2e16, 16'h2e03, 16'h2df0, 16'h2ddd, 16'h2dca, 16'h2db7, 16'h2da4, 16'h2d91, 16'h2d7e, 16'h2d6b, 16'h2d58, 16'h2d45, 16'h2d32, 16'h2d1f, 16'h2d0c, 16'h2cf9, 16'h2ce6, 16'h2cd3, 16'h2cc0, 16'h2cad, 16'h2c9a, 16'h2c87, 16'h2c74, 16'h2c61, 16'h2c4e, 16'h2c3b, 16'h2c28, 16'h2c15, 16'h2c02, 16'h2bef, 16'h2bdc, 16'h2bc9, 16'h2bb6, 16'h2ba3, 16'h2b90, 16'h2b7d, 16'h2b6a, 16'h2b57, 16'h2b44, 16'h2b31, 16'h2b1e, 16'h2b0b},
                                 {16'h2af8, 16'h2ae5, 16'h2ad2, 16'h2abf, 16'h2aac, 16'h2a99, 16'h2a86, 16'h2a73, 16'h2a60, 16'h2a4d, 16'h2a3a, 16'h2a27, 16'h2a14, 16'h2a01, 16'h29ee, 16'h29db, 16'h29c8, 16'h29b5, 16'h29a2, 16'h298f, 16'h297c, 16'h2969, 16'h2956, 16'h2943, 16'h2930, 16'h291d, 16'h290a, 16'h28f7, 16'h28e4, 16'h28e4, 16'h28e4, 16'h28ef, 16'h28fd, 16'h290b, 16'h2919, 16'h2927, 16'h2935, 16'h2943, 16'h2951, 16'h295f, 16'h296d, 16'h297b, 16'h2989, 16'h2997, 16'h29a5, 16'h29b3, 16'h29c1, 16'h29cf, 16'h29dd, 16'h29eb, 16'h29f9, 16'h2a07, 16'h2a15, 16'h2a23, 16'h2a31, 16'h2a3f, 16'h2a4d, 16'h2a5b, 16'h2a69, 16'h2a77, 16'h2a85, 16'h2a93, 16'h2aa1, 16'h2aaf},
                                 {16'h2abd, 16'h2acb, 16'h2ad9, 16'h2ae7, 16'h2af5, 16'h2b03, 16'h2b11, 16'h2b1f, 16'h2b2d, 16'h2b3b, 16'h2b49, 16'h2b57, 16'h2b65, 16'h2b73, 16'h2b81, 16'h2b8f, 16'h2b9d, 16'h2bab, 16'h2bb9, 16'h2bc7, 16'h2bd5, 16'h2be3, 16'h2bf1, 16'h2bff, 16'h2c0d, 16'h2c1b, 16'h2c29, 16'h2c37, 16'h2c45, 16'h2c53, 16'h2c61, 16'h2c6f, 16'h2c7d, 16'h2c8b, 16'h2c99, 16'h2ca7, 16'h2cb5, 16'h2cc3, 16'h2cd1, 16'h2cdf, 16'h2ced, 16'h2cfb, 16'h2d09, 16'h2d17, 16'h2d25, 16'h2d33, 16'h2d41, 16'h2d4f, 16'h2d5d, 16'h2d6b, 16'h2d79, 16'h2d87, 16'h2d95, 16'h2da3, 16'h2db1, 16'h2dbf, 16'h2dcd, 16'h2ddb, 16'h2de9, 16'h2df7, 16'h2e05, 16'h2e13, 16'h2e21, 16'h2e2f},
                                 {16'h2e3d, 16'h2e4b, 16'h2e59, 16'h2e67, 16'h2e75, 16'h2e83, 16'h2e91, 16'h2e9f, 16'h2ead, 16'h2ebb, 16'h2ec9, 16'h2ed7, 16'h2ee5, 16'h2ef3, 16'h2f01, 16'h2f0f, 16'h2f1d, 16'h2f2b, 16'h2f39, 16'h2f47, 16'h2f55, 16'h2f63, 16'h2f71, 16'h2f7f, 16'h2f8d, 16'h2f9b, 16'h2fa9, 16'h2fb7, 16'h2fc5, 16'h2fd3, 16'h2fe1, 16'h2fef, 16'h2ffd, 16'h300b, 16'h3019, 16'h3027, 16'h3035, 16'h3043, 16'h3051, 16'h305f, 16'h306d, 16'h307b, 16'h3089, 16'h3097, 16'h30a5, 16'h30b3, 16'h30c1, 16'h30cf, 16'h30dd, 16'h30eb, 16'h30f9, 16'h3107, 16'h3115, 16'h3123, 16'h3131, 16'h313f, 16'h314d, 16'h315b, 16'h3169, 16'h3177, 16'h3185, 16'h3193, 16'h31a1, 16'h31af},
                                 {16'h31bd, 16'h31cb, 16'h31d9, 16'h31e7, 16'h31f5, 16'h3203, 16'h3211, 16'h321f, 16'h322d, 16'h323b, 16'h3249, 16'h3257, 16'h3265, 16'h3273, 16'h3281, 16'h328f, 16'h329d, 16'h32ab, 16'h32b9, 16'h32c7, 16'h32d5, 16'h32e3, 16'h32f1, 16'h32ff, 16'h330d, 16'h331b, 16'h3329, 16'h3337, 16'h3345, 16'h3353, 16'h3361, 16'h336f, 16'h337d, 16'h338b, 16'h3399, 16'h33a7, 16'h33b5, 16'h33c3, 16'h33d1, 16'h33df, 16'h33ed, 16'h33fb, 16'h3409, 16'h3417, 16'h3425, 16'h3433, 16'h3441, 16'h344f, 16'h345d, 16'h346b, 16'h3479, 16'h3487, 16'h3495, 16'h34a3, 16'h34b1, 16'h34bf, 16'h34cd, 16'h34db, 16'h34e9, 16'h34f7, 16'h3505, 16'h3513, 16'h3521, 16'h352f},
                                 {16'h353d, 16'h354b, 16'h3559, 16'h3567, 16'h3575, 16'h3583, 16'h3591, 16'h359f, 16'h35ad, 16'h35bb, 16'h35c9, 16'h35d7, 16'h35e5, 16'h35f3, 16'h3601, 16'h360f, 16'h361d, 16'h362b, 16'h3639, 16'h3647, 16'h3655, 16'h3663, 16'h3671, 16'h367f, 16'h368d, 16'h369b, 16'h36a9, 16'h36b7, 16'h36c5, 16'h36d3, 16'h36e1, 16'h36ef, 16'h36fd, 16'h370b, 16'h3719, 16'h3727, 16'h3735, 16'h3743, 16'h3751, 16'h375f, 16'h376d, 16'h377b, 16'h3789, 16'h3797, 16'h37a5, 16'h37d2, 16'h37d5, 16'h37d8, 16'h37db, 16'h37de, 16'h37e1, 16'h37e4, 16'h37e7, 16'h37ea, 16'h37ed, 16'h37f0, 16'h37f3, 16'h37f6, 16'h37f9, 16'h37fc, 16'h37ff, 16'h3802, 16'h3805, 16'h3808},
                                 {16'h380b, 16'h380e, 16'h3811, 16'h3814, 16'h3817, 16'h381a, 16'h381d, 16'h3820, 16'h3823, 16'h3826, 16'h3829, 16'h382c, 16'h382f, 16'h3832, 16'h3835, 16'h3838, 16'h383b, 16'h383e, 16'h3841, 16'h3844, 16'h3847, 16'h384a, 16'h384d, 16'h3850, 16'h3853, 16'h3856, 16'h3859, 16'h385c, 16'h385f, 16'h3862, 16'h3865, 16'h3868, 16'h386b, 16'h386e, 16'h3871, 16'h3874, 16'h3877, 16'h387a, 16'h387d, 16'h3880, 16'h3883, 16'h3886, 16'h3889, 16'h388c, 16'h388f, 16'h3892, 16'h3895, 16'h3898, 16'h389b, 16'h389e, 16'h38a1, 16'h38a4, 16'h38a7, 16'h38aa, 16'h38ad, 16'h38b0, 16'h38b3, 16'h38b6, 16'h38b9, 16'h38bc, 16'h38bf, 16'h38c2, 16'h38c5, 16'h38c8},
                                 {16'h38cb, 16'h38ce, 16'h38d1, 16'h38d4, 16'h38d7, 16'h38da, 16'h38dd, 16'h38e0, 16'h38e3, 16'h38e6, 16'h38e9, 16'h38ec, 16'h38ef, 16'h38f2, 16'h38f5, 16'h38f8, 16'h38fb, 16'h38fe, 16'h3901, 16'h3904, 16'h3907, 16'h38f3, 16'h38ed, 16'h38e7, 16'h38e1, 16'h38db, 16'h38d5, 16'h38cf, 16'h38c9, 16'h38c3, 16'h38bd, 16'h38b7, 16'h38b1, 16'h38ab, 16'h38a5, 16'h389f, 16'h3899, 16'h3893, 16'h388d, 16'h3887, 16'h3881, 16'h387b, 16'h3875, 16'h386f, 16'h3869, 16'h3863, 16'h385d, 16'h3857, 16'h3851, 16'h384b, 16'h3845, 16'h383f, 16'h3839, 16'h3833, 16'h382d, 16'h3827, 16'h3821, 16'h381b, 16'h3815, 16'h380f, 16'h3809, 16'h3803, 16'h37fd, 16'h37f7},
                                 {16'h37f1, 16'h37eb, 16'h37e5, 16'h37df, 16'h37d9, 16'h37d3, 16'h37cd, 16'h37c7, 16'h37c1, 16'h37bb, 16'h37b5, 16'h37af, 16'h37a9, 16'h37a3, 16'h379d, 16'h3797, 16'h3791, 16'h378b, 16'h3785, 16'h377f, 16'h3779, 16'h3773, 16'h376d, 16'h3767, 16'h3761, 16'h375b, 16'h3755, 16'h374f, 16'h3749, 16'h3743, 16'h373d, 16'h3737, 16'h3731, 16'h372b, 16'h3725, 16'h371f, 16'h3719, 16'h3713, 16'h370d, 16'h3707, 16'h3701, 16'h36fb, 16'h36f5, 16'h36ef, 16'h36e9, 16'h36e3, 16'h36dd, 16'h36d7, 16'h36d1, 16'h36cb, 16'h36c5, 16'h36bf, 16'h36b9, 16'h36b3, 16'h36ad, 16'h36a7, 16'h36a1, 16'h369b, 16'h3695, 16'h368f, 16'h3689, 16'h3683, 16'h367d, 16'h3677},
                                 {16'h3671, 16'h366b, 16'h3665, 16'h365f, 16'h3659, 16'h3653, 16'h364d, 16'h3647, 16'h3641, 16'h363b, 16'h3635, 16'h362f, 16'h3629, 16'h3623, 16'h361d, 16'h3617, 16'h3611, 16'h360b, 16'h3605, 16'h35ff, 16'h35f9, 16'h35f3, 16'h35ed, 16'h35e7, 16'h35e1, 16'h35db, 16'h35d5, 16'h35cf, 16'h35c9, 16'h35c3, 16'h35bd, 16'h35b7, 16'h35b1, 16'h35ab, 16'h35a5, 16'h359f, 16'h3599, 16'h3593, 16'h358d, 16'h3587, 16'h3581, 16'h357b, 16'h3575, 16'h356f, 16'h3569, 16'h3563, 16'h355d, 16'h3557, 16'h3551, 16'h354b, 16'h3545, 16'h353f, 16'h35e9, 16'h35ec, 16'h35ef, 16'h35f2, 16'h35f5, 16'h35f8, 16'h35fb, 16'h35fe, 16'h3601, 16'h3604, 16'h3607, 16'h360a},
                                 {16'h360d, 16'h3610, 16'h3613, 16'h3616, 16'h3619, 16'h361c, 16'h361f, 16'h3622, 16'h3625, 16'h3628, 16'h362b, 16'h362e, 16'h3631, 16'h3634, 16'h3637, 16'h363a, 16'h363d, 16'h3640, 16'h3643, 16'h3646, 16'h3649, 16'h364c, 16'h364f, 16'h3652, 16'h3655, 16'h3658, 16'h365b, 16'h365e, 16'h3661, 16'h3664, 16'h3667, 16'h366a, 16'h366d, 16'h3670, 16'h3673, 16'h3676, 16'h3679, 16'h367c, 16'h367f, 16'h3682, 16'h3685, 16'h3688, 16'h368b, 16'h368e, 16'h3691, 16'h3694, 16'h3697, 16'h369a, 16'h369d, 16'h36a0, 16'h36a3, 16'h36a6, 16'h36a9, 16'h36ac, 16'h36af, 16'h36b2, 16'h36b5, 16'h36b8, 16'h36bb, 16'h36be, 16'h36c1, 16'h36c4, 16'h36c7, 16'h36ca},
                                 {16'h36cd, 16'h36d0, 16'h36d3, 16'h36d6, 16'h36d9, 16'h36dc, 16'h36df, 16'h36e2, 16'h36e5, 16'h36e8, 16'h36eb, 16'h36ee, 16'h36f1, 16'h36f4, 16'h36f7, 16'h36fa, 16'h36fd, 16'h3700, 16'h3703, 16'h3706, 16'h3709, 16'h370c, 16'h370f, 16'h3712, 16'h3715, 16'h3718, 16'h371b, 16'h371e, 16'h3721, 16'h3724, 16'h3727, 16'h372a, 16'h372d, 16'h3730, 16'h3733, 16'h3736, 16'h3739, 16'h373c, 16'h373f, 16'h3742, 16'h3745, 16'h3748, 16'h374b, 16'h374e, 16'h3751, 16'h3754, 16'h3757, 16'h375a, 16'h375d, 16'h3760, 16'h3763, 16'h3766, 16'h3769, 16'h376c, 16'h376f, 16'h3772, 16'h3775, 16'h3778, 16'h377b, 16'h377e, 16'h3781, 16'h3784, 16'h3787, 16'h378a},
                                 {16'h378d, 16'h3790, 16'h3793, 16'h3796, 16'h3799, 16'h379c, 16'h379f, 16'h37a2, 16'h37a5, 16'h37a8, 16'h37ab, 16'h37ae, 16'h37b1, 16'h37b4, 16'h37b7, 16'h37ba, 16'h37bd, 16'h37c0, 16'h37c3, 16'h37c6, 16'h37c9, 16'h37cc, 16'h37cf, 16'h37d2, 16'h37d5, 16'h37d8, 16'h37db, 16'h37de, 16'h37e1, 16'h37e4, 16'h37e7, 16'h37ea, 16'h37ed, 16'h37f0, 16'h37f3, 16'h37f6, 16'h37f9, 16'h37fc, 16'h37ff, 16'h3802, 16'h3805, 16'h3808, 16'h380b, 16'h380e, 16'h3811, 16'h3814, 16'h3817, 16'h381a, 16'h381d, 16'h3820, 16'h3823, 16'h3826, 16'h3829, 16'h382c, 16'h382f, 16'h3832, 16'h3835, 16'h3838, 16'h383b, 16'h383e, 16'h3841, 16'h3844, 16'h3847, 16'h384a},
                                 {16'h384d, 16'h3850, 16'h3853, 16'h3856, 16'h3859, 16'h385c, 16'h385f, 16'h3862, 16'h3865, 16'h3868, 16'h386b, 16'h386e, 16'h3871, 16'h3874, 16'h3877, 16'h387a, 16'h387d, 16'h3880, 16'h3883, 16'h3886, 16'h3889, 16'h388c, 16'h388f, 16'h3892, 16'h3895, 16'h3898, 16'h389b, 16'h389e, 16'h38a1, 16'h38a4, 16'h38a7, 16'h38aa, 16'h38ad, 16'h38b0, 16'h38b3, 16'h38b6, 16'h38b9, 16'h38bc, 16'h38bf, 16'h38c2, 16'h38c5, 16'h38c8, 16'h38cb, 16'h38ce, 16'h38d1, 16'h38d4, 16'h38d7, 16'h38da, 16'h38dd, 16'h38e0, 16'h38e3, 16'h38e6, 16'h38e9, 16'h38ec, 16'h38ef, 16'h38f2, 16'h38f5, 16'h38f8, 16'h38fb, 16'h38fe, 16'h3901, 16'h3904, 16'h3907, 16'h390a},
                                 {16'h390d, 16'h3910, 16'h3913, 16'h3916, 16'h3919, 16'h391c, 16'h391f, 16'h3922, 16'h3925, 16'h3928, 16'h392b, 16'h392e, 16'h3931, 16'h3934, 16'h3937, 16'h393a, 16'h393d, 16'h3940, 16'h3943, 16'h3946, 16'h3949, 16'h394c, 16'h394f, 16'h3952, 16'h3955, 16'h3958, 16'h395b, 16'h395e, 16'h3961, 16'h3964, 16'h3967, 16'h396a, 16'h396d, 16'h3970, 16'h3973, 16'h3976, 16'h3979, 16'h397c, 16'h397f, 16'h3982, 16'h3985, 16'h3988, 16'h398b, 16'h398e, 16'h3991, 16'h3994, 16'h3997, 16'h399a, 16'h399d, 16'h39a0, 16'h39a3, 16'h39a6, 16'h39a9, 16'h39ac, 16'h39af, 16'h39b2, 16'h39b5, 16'h39b8, 16'h39bb, 16'h39be, 16'h39c1, 16'h39c4, 16'h39c7, 16'h39ca},
                                 {16'h39cd, 16'h39d0, 16'h39d3, 16'h39d6, 16'h39d9, 16'h39dc, 16'h39df, 16'h39e2, 16'h39e5, 16'h39e8, 16'h39eb, 16'h39ee, 16'h39f1, 16'h39f4, 16'h39f7, 16'h39fa, 16'h39fd, 16'h3a00, 16'h3a03, 16'h3a06, 16'h3a09, 16'h3a0c, 16'h3a0f, 16'h3a12, 16'h3a15, 16'h3a18, 16'h3a1b, 16'h3a1e, 16'h3a21, 16'h3a24, 16'h3a27, 16'h3a2a, 16'h3a2d, 16'h3a30, 16'h3a33, 16'h3a36, 16'h3a39, 16'h3a3c, 16'h3a3f, 16'h3a42, 16'h3a45, 16'h3a48, 16'h3a4b, 16'h3a4e, 16'h3a51, 16'h3a54, 16'h3a57, 16'h3a5a, 16'h3a5d, 16'h3a60, 16'h3a63, 16'h3a66, 16'h3a69, 16'h3a6c, 16'h3a6f, 16'h3a72, 16'h3a75, 16'h3a78, 16'h3a7b, 16'h3a7e, 16'h3a6c, 16'h3a54, 16'h3a3c, 16'h3a24},
                                 {16'h3a0c, 16'h39f4, 16'h39dc, 16'h39c4, 16'h39ac, 16'h3994, 16'h397c, 16'h3964, 16'h394c, 16'h3934, 16'h391c, 16'h3904, 16'h38ec, 16'h38d4, 16'h38bc, 16'h38a4, 16'h388c, 16'h3874, 16'h385c, 16'h3844, 16'h382c, 16'h3814, 16'h37fc, 16'h37e4, 16'h37cc, 16'h37b4, 16'h379c, 16'h3784, 16'h376c, 16'h3754, 16'h373c, 16'h3724, 16'h370c, 16'h36f4, 16'h36dc, 16'h36c4, 16'h36ac, 16'h3694, 16'h367c, 16'h3664, 16'h364c, 16'h3634, 16'h361c, 16'h3604, 16'h35ec, 16'h35d4, 16'h35bc, 16'h35a4, 16'h358c, 16'h3574, 16'h355c, 16'h3544, 16'h352c, 16'h3514, 16'h34fc, 16'h34e4, 16'h34cc, 16'h34b4, 16'h349c, 16'h3484, 16'h346c, 16'h3454, 16'h343c, 16'h3424},
                                 {16'h340c, 16'h33f4, 16'h33dc, 16'h33c4, 16'h33ac, 16'h3394, 16'h337c, 16'h3364, 16'h334c, 16'h3334, 16'h331c, 16'h3304, 16'h32ec, 16'h32d4, 16'h32bc, 16'h32a4, 16'h328c, 16'h3274, 16'h325c, 16'h3244, 16'h322c, 16'h3214, 16'h31fc, 16'h31e4, 16'h31cc, 16'h31b4, 16'h319c, 16'h3184, 16'h316c, 16'h3154, 16'h313c, 16'h3124, 16'h310c, 16'h30f4, 16'h30dc, 16'h30c4, 16'h30ac, 16'h3094, 16'h307c, 16'h3064, 16'h304c, 16'h3034, 16'h301c, 16'h3004, 16'h2fec, 16'h2fd4, 16'h2fbc, 16'h2fa4, 16'h2f8c, 16'h2f74, 16'h2f5c, 16'h2f44, 16'h2f2c, 16'h2f14, 16'h2efc, 16'h2ee4, 16'h2ecc, 16'h2eb4, 16'h2e9c, 16'h2e84, 16'h2e6c, 16'h2e54, 16'h2e3c, 16'h2e24},
                                 {16'h2e0c, 16'h2df4, 16'h2ddc, 16'h2dc4, 16'h2dac, 16'h2d94, 16'h2d7c, 16'h2d64, 16'h2d4c, 16'h2d34, 16'h2d1c, 16'h2d04, 16'h2cec, 16'h2cd4, 16'h2cbc, 16'h2ca4, 16'h2c8c, 16'h2c74, 16'h2c5c, 16'h2c44, 16'h2c2c, 16'h2c14, 16'h2bfc, 16'h2be4, 16'h2bcc, 16'h2bb4, 16'h2b9c, 16'h2b84, 16'h2b6c, 16'h2b54, 16'h2b3c, 16'h2b24, 16'h2b0c, 16'h2af4, 16'h2adc, 16'h2ac4, 16'h2aac, 16'h2a94, 16'h2a7c, 16'h2a64, 16'h2a4c, 16'h2a34, 16'h2a1c, 16'h2a04, 16'h29ec, 16'h29d4, 16'h29bc, 16'h29a4, 16'h298c, 16'h2974, 16'h295c, 16'h2944, 16'h292c, 16'h2914, 16'h28fc, 16'h28e4, 16'h28cc, 16'h28b4, 16'h289c, 16'h2884, 16'h286c, 16'h2854, 16'h283c, 16'h2824},
                                 {16'h280c, 16'h27f4, 16'h27dc, 16'h27c4, 16'h27ac, 16'h2794, 16'h277c, 16'h2764, 16'h274c, 16'h2734, 16'h271c, 16'h2704, 16'h26ec, 16'h26d4, 16'h26bc, 16'h26a4, 16'h268c, 16'h2674, 16'h265c, 16'h2644, 16'h262c, 16'h2614, 16'h25fc, 16'h25e4, 16'h25cc, 16'h25b4, 16'h259c, 16'h2584, 16'h256c, 16'h2554, 16'h253c, 16'h2524, 16'h250c, 16'h24f4, 16'h24dc, 16'h24c4, 16'h24ac, 16'h2494, 16'h247c, 16'h2464, 16'h244c, 16'h2434, 16'h241c, 16'h2404, 16'h23ec, 16'h23d4, 16'h23bc, 16'h23a4, 16'h238c, 16'h2374, 16'h235c, 16'h2344, 16'h232c, 16'h2314, 16'h22fc, 16'h22e4, 16'h22cc, 16'h22b4, 16'h229c, 16'h2284, 16'h226c, 16'h2254, 16'h223c, 16'h2224},
                                 {16'h220c, 16'h21f4, 16'h21dc, 16'h21c4, 16'h21ac, 16'h2194, 16'h217c, 16'h2164, 16'h214c, 16'h2134, 16'h211c, 16'h2104, 16'h20ec, 16'h20d4, 16'h20bc, 16'h20a4, 16'h208c, 16'h2074, 16'h205c, 16'h2044, 16'h202c, 16'h2014, 16'h1ffc, 16'h1fe4, 16'h1fcc, 16'h1fb4, 16'h1f9c, 16'h1f84, 16'h1f6c, 16'h1f54, 16'h1f3c, 16'h1f24, 16'h1f0c, 16'h1ef4, 16'h1edc, 16'h1ec4, 16'h1eac, 16'h1e94, 16'h1e7c, 16'h1e64, 16'h1e4c, 16'h1e34, 16'h1e1c, 16'h1e04, 16'h1dec, 16'h1dd4, 16'h1dbc, 16'h1da4, 16'h1d8c, 16'h1d74, 16'h1d5c, 16'h1d44, 16'h1d2c, 16'h1d14, 16'h1cfc, 16'h1ce4, 16'h1ccc, 16'h1cb4, 16'h1c9c, 16'h1ce4, 16'h1d1d, 16'h1d56, 16'h1d8f, 16'h1dc8},
                                 {16'h1e01, 16'h1e3a, 16'h1e73, 16'h1eac, 16'h1ee5, 16'h1f1e, 16'h1f57, 16'h1f90, 16'h1fc9, 16'h2002, 16'h203b, 16'h2074, 16'h20ad, 16'h20e6, 16'h211f, 16'h2158, 16'h2191, 16'h21ca, 16'h2203, 16'h223c, 16'h2275, 16'h22ae, 16'h22e7, 16'h2320, 16'h2359, 16'h2392, 16'h23cb, 16'h2404, 16'h243d, 16'h2476, 16'h24af, 16'h24e8, 16'h2521, 16'h255a, 16'h2593, 16'h2593, 16'h2597, 16'h259f, 16'h25a7, 16'h25af, 16'h25b7, 16'h25bf, 16'h25c7, 16'h25cf, 16'h25d7, 16'h25df, 16'h25e7, 16'h25ef, 16'h25f7, 16'h25ff, 16'h2607, 16'h260f, 16'h2617, 16'h261f, 16'h2627, 16'h262f, 16'h2637, 16'h263f, 16'h2647, 16'h264f, 16'h2657, 16'h265f, 16'h2667, 16'h266f},
                                 {16'h2677, 16'h267f, 16'h2687, 16'h268f, 16'h2697, 16'h269f, 16'h26a7, 16'h26af, 16'h26b7, 16'h26bf, 16'h26c7, 16'h26cf, 16'h26d7, 16'h26df, 16'h26e7, 16'h26ef, 16'h26f7, 16'h26ff, 16'h2707, 16'h270f, 16'h2717, 16'h271f, 16'h2727, 16'h272f, 16'h2737, 16'h273f, 16'h2747, 16'h274f, 16'h2757, 16'h275f, 16'h2767, 16'h276f, 16'h2777, 16'h277f, 16'h2787, 16'h278f, 16'h2797, 16'h279f, 16'h27a7, 16'h27af, 16'h27b7, 16'h27bf, 16'h27c7, 16'h27cf, 16'h27d7, 16'h27df, 16'h27e7, 16'h27ef, 16'h27f7, 16'h27ff, 16'h2807, 16'h280f, 16'h2817, 16'h281f, 16'h2827, 16'h282f, 16'h2837, 16'h283f, 16'h2847, 16'h284f, 16'h2857, 16'h285f, 16'h2867, 16'h286f},
                                 {16'h2877, 16'h287f, 16'h2887, 16'h288f, 16'h2897, 16'h289f, 16'h28a7, 16'h28af, 16'h28b7, 16'h28bf, 16'h28c7, 16'h28cf, 16'h28d7, 16'h28df, 16'h28e7, 16'h28ef, 16'h28f7, 16'h28ff, 16'h2907, 16'h290f, 16'h2917, 16'h291f, 16'h2927, 16'h292f, 16'h2937, 16'h293f, 16'h2947, 16'h294f, 16'h2957, 16'h295f, 16'h2967, 16'h296f, 16'h2977, 16'h297f, 16'h2987, 16'h298f, 16'h2997, 16'h299f, 16'h29a7, 16'h29af, 16'h29b7, 16'h29bf, 16'h29c7, 16'h29cf, 16'h29d7, 16'h29df, 16'h29e7, 16'h29ef, 16'h29f7, 16'h29ff, 16'h2a07, 16'h2a0f, 16'h2a17, 16'h2a1f, 16'h2a27, 16'h2a2f, 16'h2a37, 16'h2a3f, 16'h2a47, 16'h2a4f, 16'h2a57, 16'h2a5f, 16'h2a67, 16'h2a6f},
                                 {16'h2a77, 16'h2a7f, 16'h2a87, 16'h2a8f, 16'h2a97, 16'h2a9f, 16'h2aa7, 16'h2aaf, 16'h2ab7, 16'h2abf, 16'h2ac7, 16'h2acf, 16'h2ad7, 16'h2adf, 16'h2ae7, 16'h2aef, 16'h2af7, 16'h2aff, 16'h2b07, 16'h2b0f, 16'h2b17, 16'h2b1f, 16'h2b27, 16'h2b2f, 16'h2b37, 16'h2b3f, 16'h2b47, 16'h2b4f, 16'h2b57, 16'h2b5f, 16'h2b67, 16'h2b6f, 16'h2b77, 16'h2b7f, 16'h2b87, 16'h2b8f, 16'h2b97, 16'h2b9f, 16'h2ba7, 16'h2baf, 16'h2bb7, 16'h2bbf, 16'h2bc7, 16'h2bcf, 16'h2bd7, 16'h2bdf, 16'h2be7, 16'h2bef, 16'h2bf7, 16'h2bff, 16'h2c07, 16'h2c0f, 16'h2c17, 16'h2c1f, 16'h2c27, 16'h2c2f, 16'h2c37, 16'h2c3f, 16'h2c47, 16'h2c4f, 16'h2c57, 16'h2c5f, 16'h2c67, 16'h2c6f},
                                 {16'h2c77, 16'h2c7f, 16'h2c87, 16'h2c8f, 16'h2c97, 16'h2c9f, 16'h2ca7, 16'h2caf, 16'h2cb7, 16'h2cbf, 16'h2cc7, 16'h2ccf, 16'h2cd7, 16'h2cdf, 16'h2ce7, 16'h2cef, 16'h2cf7, 16'h2cff, 16'h2d07, 16'h2d0f, 16'h2d17, 16'h2d1f, 16'h2d27, 16'h2d2f, 16'h2d37, 16'h2d3f, 16'h2d47, 16'h2d4f, 16'h2d57, 16'h2d5f, 16'h2d67, 16'h2d6f, 16'h2d77, 16'h2d7f, 16'h2d7f, 16'h2d7f, 16'h2d7f, 16'h2d7f, 16'h2d7f, 16'h2d7f, 16'h2d7a, 16'h2d69, 16'h2d58, 16'h2d47, 16'h2d36, 16'h2d25, 16'h2d14, 16'h2d03, 16'h2cf2, 16'h2ce1, 16'h2cd0, 16'h2cbf, 16'h2cae, 16'h2c9d, 16'h2c8c, 16'h2c7b, 16'h2c6a, 16'h2c59, 16'h2c48, 16'h2c37, 16'h2c26, 16'h2c15, 16'h2c04, 16'h2bf3},
                                 {16'h2be2, 16'h2bd1, 16'h2bc0, 16'h2baf, 16'h2b9e, 16'h2b8d, 16'h2b7c, 16'h2b6b, 16'h2b5a, 16'h2b49, 16'h2b38, 16'h2b27, 16'h2b16, 16'h2b05, 16'h2af4, 16'h2ae3, 16'h2ad2, 16'h2ac1, 16'h2ab0, 16'h2a9f, 16'h2a8e, 16'h2a7d, 16'h2a6c, 16'h2a5b, 16'h2a4a, 16'h2a39, 16'h2a28, 16'h2a17, 16'h2a06, 16'h29f5, 16'h29e4, 16'h29d3, 16'h29c2, 16'h29b1, 16'h29a0, 16'h298f, 16'h297e, 16'h296d, 16'h295c, 16'h294b, 16'h293a, 16'h2929, 16'h2918, 16'h2907, 16'h28f6, 16'h28e5, 16'h28d4, 16'h28c3, 16'h28b2, 16'h28a1, 16'h2890, 16'h287f, 16'h286e, 16'h285d, 16'h284c, 16'h283b, 16'h282a, 16'h2819, 16'h2808, 16'h27f7, 16'h27e6, 16'h27d5, 16'h27c4, 16'h27b3},
                                 {16'h27a2, 16'h2791, 16'h2780, 16'h276f, 16'h275e, 16'h274d, 16'h273c, 16'h272b, 16'h271a, 16'h2709, 16'h26f8, 16'h26e7, 16'h26d6, 16'h26c5, 16'h26b4, 16'h26a3, 16'h2692, 16'h2681, 16'h2670, 16'h265f, 16'h264e, 16'h263d, 16'h262c, 16'h261b, 16'h260a, 16'h25f9, 16'h25e8, 16'h25d7, 16'h25c6, 16'h25b5, 16'h25a4, 16'h2593, 16'h2582, 16'h2571, 16'h2560, 16'h254f, 16'h253e, 16'h252d, 16'h251c, 16'h250b, 16'h24fa, 16'h24e9, 16'h24d8, 16'h24c7, 16'h24b6, 16'h24a5, 16'h2494, 16'h2483, 16'h2472, 16'h2461, 16'h2450, 16'h243f, 16'h242e, 16'h241d, 16'h240c, 16'h23fb, 16'h23ea, 16'h23d9, 16'h23c8, 16'h23b7, 16'h23a6, 16'h2395, 16'h2384, 16'h2373},
                                 {16'h2362, 16'h2351, 16'h2340, 16'h232f, 16'h231e, 16'h230d, 16'h22fc, 16'h22eb, 16'h22da, 16'h22c9, 16'h22b8, 16'h22a7, 16'h2296, 16'h2285, 16'h2274, 16'h2263, 16'h2252, 16'h2241, 16'h2230, 16'h221f, 16'h220e, 16'h21fd, 16'h21ec, 16'h21db, 16'h21ca, 16'h21b9, 16'h21a8, 16'h2197, 16'h2186, 16'h2175, 16'h2164, 16'h2153, 16'h2142, 16'h2131, 16'h2120, 16'h210f, 16'h20fe, 16'h20ed, 16'h20dc, 16'h20cb, 16'h20ba, 16'h20a9, 16'h2098, 16'h2087, 16'h2076, 16'h2065, 16'h2054, 16'h2043, 16'h2032, 16'h2021, 16'h2010, 16'h1fff, 16'h1fee, 16'h1fdd, 16'h1fcc, 16'h1fbb, 16'h1faa, 16'h1f99, 16'h1f88, 16'h1f77, 16'h1f66, 16'h1f55, 16'h1f44, 16'h1f33},
                                 {16'h1f22, 16'h1f11, 16'h1f00, 16'h1eef, 16'h1ede, 16'h1ecd, 16'h1ebc, 16'h1eab, 16'h1e9a, 16'h1e89, 16'h1e78, 16'h1e67, 16'h1e56, 16'h1e45, 16'h1e34, 16'h1e23, 16'h1e12, 16'h1e01, 16'h1df0, 16'h1ddf, 16'h1dce, 16'h1dbd, 16'h1dac, 16'h1d9b, 16'h1d8a, 16'h1d79, 16'h1d68, 16'h1d57, 16'h1d46, 16'h1d35, 16'h1d24, 16'h1d13, 16'h1d02, 16'h1cf1, 16'h1ce0, 16'h1ccf, 16'h1cbe, 16'h1cad, 16'h1c9c, 16'h1c8b, 16'h1c7a, 16'h1c69, 16'h1c58, 16'h1c47, 16'h1c36, 16'h1c25, 16'h1c14, 16'h1c03, 16'h1bf2, 16'h1be1, 16'h1bd0, 16'h1bbf, 16'h1bae, 16'h1b9d, 16'h1b8c, 16'h1b7b, 16'h1b6a, 16'h1b59, 16'h1b48, 16'h1b37, 16'h1b26, 16'h1b15, 16'h1b04, 16'h1af3},
                                 {16'h1ae2, 16'h1ad1, 16'h1ac0, 16'h1aaf, 16'h1a9e, 16'h1a8d, 16'h1a7c, 16'h1a6b, 16'h1a5a, 16'h1a49, 16'h1a38, 16'h1a27, 16'h1a16, 16'h1a05, 16'h19f4, 16'h19e3, 16'h19d2, 16'h19c1, 16'h19b0, 16'h199f, 16'h198e, 16'h197d, 16'h196c, 16'h195b, 16'h194a, 16'h1939, 16'h1928, 16'h1917, 16'h1906, 16'h18f5, 16'h18e4, 16'h18d3, 16'h18c2, 16'h18b1, 16'h18a0, 16'h188f, 16'h187e, 16'h186d, 16'h185c, 16'h184b, 16'h183a, 16'h1829, 16'h1818, 16'h1807, 16'h17f6, 16'h17e5, 16'h17d4, 16'h17c3, 16'h17b2, 16'h17a1, 16'h1790, 16'h177f, 16'h176e, 16'h175d, 16'h174c, 16'h173b, 16'h172a, 16'h1719, 16'h1708, 16'h16f7, 16'h16e6, 16'h16d5, 16'h16c4, 16'h16b3},
                                 {16'h16a2, 16'h1691, 16'h1680, 16'h166f, 16'h165e, 16'h164d, 16'h163c, 16'h162b, 16'h161a, 16'h1609, 16'h15f8, 16'h15e7, 16'h15d6, 16'h15c5, 16'h15b4, 16'h15a3, 16'h1592, 16'h1581, 16'h1570, 16'h155f, 16'h154e, 16'h153d, 16'h152c, 16'h151b, 16'h150a, 16'h14f9, 16'h14e8, 16'h14d7, 16'h14c6, 16'h14b5, 16'h14a4, 16'h1493, 16'h1482, 16'h1471, 16'h1460, 16'h144f, 16'h143e, 16'h142d, 16'h141c, 16'h140b, 16'h13fa, 16'h13e9, 16'h13d8, 16'h13c7, 16'h13b6, 16'h13a5, 16'h1394, 16'h1383, 16'h1372, 16'h1361, 16'h1350, 16'h133f, 16'h132e, 16'h131d, 16'h130c, 16'h12fb, 16'h12ea, 16'h12d9, 16'h12c8, 16'h12b7, 16'h12a6, 16'h1295, 16'h1284, 16'h1273},
                                 {16'h1262, 16'h1251, 16'h1240, 16'h122f, 16'h121e, 16'h120d, 16'h11fc, 16'h11eb, 16'h11da, 16'h11c9, 16'h11b8, 16'h11a7, 16'h1196, 16'h1185, 16'h1174, 16'h1163, 16'h1152, 16'h1141, 16'h1130, 16'h111f, 16'h110e, 16'h10fd, 16'h10ec, 16'h10db, 16'h10ca, 16'h10b9, 16'h10a8, 16'h1097, 16'h1086, 16'h1075, 16'h1064, 16'h1053, 16'h1042, 16'h1031, 16'h1020, 16'h100f, 16'h0ffe, 16'h0fed, 16'h0fdc, 16'h0fcb, 16'h0fba, 16'h0fa9, 16'h0f98, 16'h0f87, 16'h0f76, 16'h0f65, 16'h0f54, 16'h0f43, 16'h0f32, 16'h0f21, 16'h0f10, 16'h0eff, 16'h0eee, 16'h0edd, 16'h0ecc, 16'h0ebb, 16'h0eaa, 16'h0e99, 16'h0e88, 16'h0e77, 16'h0e66, 16'h0e55, 16'h0e44, 16'h0e33},
                                 {16'h0e22, 16'h0e11, 16'h0e00, 16'h0def, 16'h0dde, 16'h0dcd, 16'h0dbc, 16'h0dab, 16'h0d9a, 16'h0d89, 16'h0d78, 16'h0d67, 16'h0d56, 16'h0d45, 16'h0d34, 16'h0d23, 16'h0d12, 16'h0d01, 16'h0cf0, 16'h0cdf, 16'h0cce, 16'h0cbd, 16'h0cac, 16'h0c9b, 16'h0c8a, 16'h0c79, 16'h0c68, 16'h0c57, 16'h0c46, 16'h0c35, 16'h0c24, 16'h0c13, 16'h0c02, 16'h0bf1, 16'h0be0, 16'h0bcf, 16'h0bbe, 16'h0bad, 16'h0b9c, 16'h0b8b, 16'h0b7a, 16'h0b69, 16'h0b58, 16'h0b47, 16'h0b36, 16'h0b25, 16'h0b14, 16'h0b03, 16'h0af2, 16'h0ae1, 16'h0ad0, 16'h0abf, 16'h0aae, 16'h0a9d, 16'h0a8c, 16'h0a7b, 16'h0a6a, 16'h0a59, 16'h0a48, 16'h0a37, 16'h0a26, 16'h0a15, 16'h0a04, 16'h09f3},
                                 {16'h09e2, 16'h09d1, 16'h09c0, 16'h09af, 16'h099e, 16'h098d, 16'h097c, 16'h096b, 16'h095a, 16'h0949, 16'h0938, 16'h0927, 16'h0916, 16'h0905, 16'h08f4, 16'h08e3, 16'h08d2, 16'h08c1, 16'h08b0, 16'h089f, 16'h088e, 16'h087d, 16'h086c, 16'h085b, 16'h084a, 16'h0839, 16'h0828, 16'h0817, 16'h0806, 16'h07f5, 16'h07e4, 16'h07d3, 16'h07c2, 16'h07b1, 16'h07a0, 16'h078f, 16'h077e, 16'h076d, 16'h075c, 16'h074b, 16'h073a, 16'h0729, 16'h0718, 16'h0707, 16'h06f6, 16'h06e5, 16'h06d4, 16'h06c3, 16'h06b2, 16'h06a1, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690},
                                 {16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690},
                                 {16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690},
                                 {16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h0690, 16'h068f},
                                 {16'h068e, 16'h068d, 16'h068c, 16'h068b, 16'h068a, 16'h0689, 16'h0688, 16'h0687, 16'h0686, 16'h0685, 16'h0684, 16'h0683, 16'h0682, 16'h0681, 16'h0680, 16'h067f, 16'h067e, 16'h067d, 16'h067c, 16'h067b, 16'h067a, 16'h0679, 16'h0678, 16'h0677, 16'h0676, 16'h0675, 16'h0674, 16'h0673, 16'h0672, 16'h0671, 16'h0670, 16'h066f, 16'h066e, 16'h066d, 16'h06aa, 16'h06c1, 16'h06d8, 16'h06ef, 16'h0706, 16'h071d, 16'h0734, 16'h074b, 16'h0762, 16'h0779, 16'h0790, 16'h07a7, 16'h07be, 16'h07d5, 16'h07ec, 16'h0803, 16'h081a, 16'h0831, 16'h0848, 16'h085f, 16'h0876, 16'h088d, 16'h08a4, 16'h08bb, 16'h08d2, 16'h08e9, 16'h0900, 16'h0917, 16'h092e, 16'h0945},
                                 {16'h095c, 16'h0973, 16'h098a, 16'h09a1, 16'h09b8, 16'h09cf, 16'h09e6, 16'h09fd, 16'h0a14, 16'h0a2b, 16'h0a42, 16'h0a59, 16'h0a70, 16'h0a87, 16'h0a9e, 16'h0ab5, 16'h0acc, 16'h0ae3, 16'h0afa, 16'h0b11, 16'h0b28, 16'h0b3f, 16'h0b56, 16'h0b6d, 16'h0b84, 16'h0b9b, 16'h0bb2, 16'h0bc9, 16'h0be0, 16'h0bf7, 16'h0c0e, 16'h0c25, 16'h0c3c, 16'h0c53, 16'h0c6a, 16'h0c81, 16'h0c98, 16'h0caf, 16'h0cc6, 16'h0cdd, 16'h0cf4, 16'h0d0b, 16'h0d22, 16'h0d39, 16'h0d50, 16'h0d67, 16'h0d7e, 16'h0d95, 16'h0dac, 16'h0dc3, 16'h0dda, 16'h0df1, 16'h0e08, 16'h0e1f, 16'h0e36, 16'h0e4d, 16'h0e64, 16'h0e7b, 16'h0e92, 16'h0ea9, 16'h0ec0, 16'h0ed7, 16'h0eee, 16'h0f05},
                                 {16'h0f1c, 16'h0f33, 16'h0f4a, 16'h0f61, 16'h0f78, 16'h0f8f, 16'h0fa6, 16'h0fbd, 16'h0fd4, 16'h0feb, 16'h1002, 16'h1019, 16'h1030, 16'h1047, 16'h105e, 16'h1075, 16'h108c, 16'h10a3, 16'h10ba, 16'h10d1, 16'h10fa, 16'h1111, 16'h1128, 16'h113f, 16'h1156, 16'h116d, 16'h1184, 16'h119b, 16'h11b2, 16'h11c9, 16'h11e0, 16'h11f7, 16'h120e, 16'h1225, 16'h123c, 16'h1253, 16'h126a, 16'h1281, 16'h1298, 16'h12af, 16'h12c6, 16'h12dd, 16'h12f4, 16'h130b, 16'h1322, 16'h1339, 16'h1350, 16'h1367, 16'h137e, 16'h1395, 16'h13ac, 16'h13c3, 16'h13da, 16'h13f1, 16'h1408, 16'h141f, 16'h1436, 16'h144d, 16'h1464, 16'h147b, 16'h1492, 16'h14a9, 16'h14c0, 16'h14d7},
                                 {16'h14ee, 16'h1505, 16'h151c, 16'h1533, 16'h154a, 16'h1561, 16'h1578, 16'h158f, 16'h15a6, 16'h15bd, 16'h15d4, 16'h15eb, 16'h1602, 16'h1619, 16'h1630, 16'h1647, 16'h165e, 16'h1675, 16'h168c, 16'h16a3, 16'h16ba, 16'h16d1, 16'h16e8, 16'h16ff, 16'h1716, 16'h172d, 16'h1744, 16'h175b, 16'h1772, 16'h1789, 16'h17a0, 16'h17b7, 16'h17ce, 16'h17e5, 16'h17fc, 16'h1813, 16'h182a, 16'h1841, 16'h1858, 16'h186f, 16'h1886, 16'h189d, 16'h18b4, 16'h18cb, 16'h18e2, 16'h18f9, 16'h1910, 16'h1927, 16'h193e, 16'h1955, 16'h196c, 16'h1983, 16'h199a, 16'h19b1, 16'h19c8, 16'h19df, 16'h19f6, 16'h1a0d, 16'h1a24, 16'h1a3b, 16'h1a52, 16'h1a69, 16'h1a80, 16'h1a97},
                                 {16'h1aae, 16'h1ac5, 16'h1adc, 16'h1af3, 16'h1b0a, 16'h1b21, 16'h1b38, 16'h1b4f, 16'h1b66, 16'h1b7d, 16'h1b94, 16'h1bab, 16'h1bc2, 16'h1bd9, 16'h1bf0, 16'h1c07, 16'h1c1e, 16'h1c35, 16'h1c4c, 16'h1c63, 16'h1c7a, 16'h1c91, 16'h1ca8, 16'h1cbf, 16'h1cd6, 16'h1ced, 16'h1d04, 16'h1d1b, 16'h1d32, 16'h1d49, 16'h1d60, 16'h1d77, 16'h1d8e, 16'h1da5, 16'h1dbc, 16'h1dd3, 16'h1dea, 16'h1e01, 16'h1e18, 16'h1e2f, 16'h1e46, 16'h1e5d, 16'h1e74, 16'h1e8b, 16'h1ea2, 16'h1eb9, 16'h1ed0, 16'h1ee7, 16'h1efe, 16'h1f15, 16'h1f2c, 16'h1f43, 16'h1f5a, 16'h1f71, 16'h1f88, 16'h1f9f, 16'h1fb6, 16'h1fcd, 16'h1fe4, 16'h1ffb, 16'h2012, 16'h2029, 16'h2040, 16'h2057},
                                 {16'h206e, 16'h2085, 16'h209c, 16'h20b3, 16'h20ca, 16'h20e1, 16'h20f8, 16'h210f, 16'h2126, 16'h213d, 16'h2154, 16'h216b, 16'h2182, 16'h2199, 16'h21b0, 16'h21c7, 16'h21de, 16'h21f5, 16'h220c, 16'h2223, 16'h223a, 16'h2251, 16'h2268, 16'h227f, 16'h2296, 16'h22ad, 16'h22c4, 16'h22db, 16'h22f2, 16'h2309, 16'h2320, 16'h2337, 16'h234e, 16'h2365, 16'h237c, 16'h2393, 16'h23aa, 16'h23c1, 16'h23d8, 16'h23ef, 16'h2406, 16'h241d, 16'h2434, 16'h244b, 16'h2462, 16'h2479, 16'h2490, 16'h24a7, 16'h24be, 16'h24d5, 16'h24ec, 16'h2503, 16'h251a, 16'h2531, 16'h2548, 16'h255f, 16'h2576, 16'h258d, 16'h25a4, 16'h25bb, 16'h25d2, 16'h25e9, 16'h2600, 16'h2617},
                                 {16'h262e, 16'h2645, 16'h265c, 16'h2673, 16'h268a, 16'h26a1, 16'h26b8, 16'h26cf, 16'h26e6, 16'h26fd, 16'h2714, 16'h272b, 16'h2742, 16'h0a32, 16'h0a32, 16'h0a32, 16'h0a32, 16'h0a32, 16'h0a32, 16'h0a32, 16'h0a32, 16'h0a32, 16'h0a32, 16'h0a32, 16'h0a32, 16'h0a32, 16'h0a32, 16'h0a32, 16'h0a32, 16'h0a2c, 16'h0a24, 16'h0a1c, 16'h0a14, 16'h0a0c, 16'h0a04, 16'h09fc, 16'h09f4, 16'h09ec, 16'h09e4, 16'h09dc, 16'h09d4, 16'h09cc, 16'h09c4, 16'h09bc, 16'h09b4, 16'h09ac, 16'h09a4, 16'h099c, 16'h0994, 16'h098c, 16'h0984, 16'h097c, 16'h0974, 16'h096c, 16'h0964, 16'h095c, 16'h0954, 16'h094c, 16'h0944, 16'h093c, 16'h0934, 16'h092c, 16'h0924, 16'h091c},
                                 {16'h0914, 16'h090c, 16'h0904, 16'h08fc, 16'h08f4, 16'h08ec, 16'h08e4, 16'h08dc, 16'h08d4, 16'h08cc, 16'h08c4, 16'h08bc, 16'h08b4, 16'h08ac, 16'h08a4, 16'h089c, 16'h0894, 16'h088c, 16'h0884, 16'h087c, 16'h0874, 16'h086c, 16'h0864, 16'h085c, 16'h0854, 16'h084c, 16'h0844, 16'h083c, 16'h0834, 16'h082c, 16'h0824, 16'h081c, 16'h0814, 16'h080c, 16'h0804, 16'h07fc, 16'h07f4, 16'h07ec, 16'h07e4, 16'h07dc, 16'h07d4, 16'h07cc, 16'h07c4, 16'h07bc, 16'h07b4, 16'h07ac, 16'h07a4, 16'h079c, 16'h0794, 16'h078c, 16'h0784, 16'h077c, 16'h0774, 16'h076c, 16'h0764, 16'h075c, 16'h0754, 16'h074c, 16'h0744, 16'h073c, 16'h0734, 16'h072c, 16'h0724, 16'h071c},
                                 {16'h0714, 16'h070c, 16'h0704, 16'h06fc, 16'h06f4, 16'h06ec, 16'h06e4, 16'h06dc, 16'h06d4, 16'h06cc, 16'h06c4, 16'h06bc, 16'h06b4, 16'h06ac, 16'h06a4, 16'h069c, 16'h0694, 16'h068c, 16'h0684, 16'h067c, 16'h0674, 16'h066c, 16'h0664, 16'h065c, 16'h0654, 16'h064c, 16'h0644, 16'h063c, 16'h0634, 16'h062c, 16'h0624, 16'h061c, 16'h0614, 16'h060c, 16'h0604, 16'h05fc, 16'h05f4, 16'h05ec, 16'h05e4, 16'h05dc, 16'h05d4, 16'h05cc, 16'h05c4, 16'h05bc, 16'h05b4, 16'h05ac, 16'h05a4, 16'h059c, 16'h0594, 16'h058c, 16'h0584, 16'h057c, 16'h0574, 16'h056c, 16'h0564, 16'h055c, 16'h0554, 16'h054c, 16'h0544, 16'h053c, 16'h0534, 16'h052c, 16'h0524, 16'h051c},
                                 {16'h0514, 16'h050c, 16'h0504, 16'h04fc, 16'h04f4, 16'h04ec, 16'h04e4, 16'h04dc, 16'h04d4, 16'h04cc, 16'h04c4, 16'h04bc, 16'h04b4, 16'h04ac, 16'h04a4, 16'h049c, 16'h0494, 16'h048c, 16'h0484, 16'h047c, 16'h0474, 16'h046c, 16'h0464, 16'h045c, 16'h0454, 16'h044c, 16'h0444, 16'h043c, 16'h0434, 16'h042c, 16'h0424, 16'h041c, 16'h0414, 16'h040c, 16'h0404, 16'h03fc, 16'h03f4, 16'h03ec, 16'h03e4, 16'h03dc, 16'h03d4, 16'h03cc, 16'h03c4, 16'h03bc, 16'h03b4, 16'h03ac, 16'h03a4, 16'h039c, 16'h0394, 16'h038c, 16'h0384, 16'h037c, 16'h0374, 16'h036c, 16'h0364, 16'h035c, 16'h0354, 16'h034c, 16'h0344, 16'h033c, 16'h0334, 16'h032c, 16'h0324, 16'h031c},
                                 {16'h0314, 16'h030c, 16'h0304, 16'h02fc, 16'h02f4, 16'h02ec, 16'h02e4, 16'h02dc, 16'h02d4, 16'h02cc, 16'h02c4, 16'h02bc, 16'h02b4, 16'h02ac, 16'h02a4, 16'h029c, 16'h0294, 16'h028c, 16'h0284, 16'h027c, 16'h0274, 16'h026c, 16'h0264, 16'h025c, 16'h0254, 16'h024c, 16'h0244, 16'h023c, 16'h0234, 16'h022c, 16'h0224, 16'h021c, 16'h0214, 16'h020c, 16'h0204, 16'h01fc, 16'h01f4, 16'h01ec, 16'h025f, 16'h029a, 16'h02d5, 16'h0310, 16'h034b, 16'h0386, 16'h03c1, 16'h03fc, 16'h0437, 16'h0472, 16'h04ad, 16'h04e8, 16'h0523, 16'h055e, 16'h0599, 16'h05d4, 16'h060f, 16'h064a, 16'h0685, 16'h06c0, 16'h06fb, 16'h0736, 16'h0771, 16'h07ac, 16'h07e7, 16'h0822},
                                 {16'h085d, 16'h0898, 16'h08d3, 16'h090e, 16'h0949, 16'h0984, 16'h09bf, 16'h09fa, 16'h0a35, 16'h0a70, 16'h0aab, 16'h0ae6, 16'h0b21, 16'h0b5c, 16'h0b97, 16'h0bd2, 16'h0c0d, 16'h0c48, 16'h0c83, 16'h0cbe, 16'h0cf9, 16'h0d34, 16'h0d6f, 16'h0daa, 16'h0de5, 16'h0e20, 16'h0e5b, 16'h0e96, 16'h0ed1, 16'h0f0c, 16'h0f47, 16'h0f82, 16'h0fbd, 16'h0ff8, 16'h1033, 16'h106e, 16'h10a9, 16'h10e4, 16'h111f, 16'h115a, 16'h1195, 16'h11d0, 16'h120b, 16'h1246, 16'h1281, 16'h12bc, 16'h12f7, 16'h1332, 16'h136d, 16'h13a8, 16'h13e3, 16'h141e, 16'h1459, 16'h1494, 16'h14cf, 16'h150a, 16'h1545, 16'h1580, 16'h15bb, 16'h15f6, 16'h1631, 16'h166c, 16'h16a7, 16'h16e2},
                                 {16'h171d, 16'h1758, 16'h1793, 16'h17ce, 16'h1809, 16'h1844, 16'h187f, 16'h18ba, 16'h18f5, 16'h1930, 16'h196b, 16'h19a6, 16'h19e1, 16'h1a1c, 16'h1a57, 16'h1a92, 16'h1acd, 16'h1b08, 16'h1b43, 16'h1b7e, 16'h1bb9, 16'h1bf4, 16'h1c2f, 16'h1c6a, 16'h1ca5, 16'h1ce0, 16'h1d1b, 16'h1d56, 16'h1d91, 16'h1dcc, 16'h1e07, 16'h1e42, 16'h1e7d, 16'h1eb8, 16'h1ef3, 16'h1f2e, 16'h1f69, 16'h1fa4, 16'h1fdf, 16'h201a, 16'h2055, 16'h2090, 16'h20cb, 16'h2106, 16'h2141, 16'h217c, 16'h21b7, 16'h21f2, 16'h222d, 16'h2268, 16'h22a3, 16'h22de, 16'h2319, 16'h2354, 16'h238f, 16'h23ca, 16'h2405, 16'h2405, 16'h2405, 16'h2405, 16'h2405, 16'h2405, 16'h2405, 16'h2405},
                                 {16'h2405, 16'h2405, 16'h2405, 16'h2405, 16'h2405, 16'h2405, 16'h2405, 16'h2405, 16'h2405, 16'h2405, 16'h2405, 16'h2401, 16'h23fc, 16'h23f7, 16'h23f2, 16'h23ed, 16'h23e8, 16'h23e3, 16'h23de, 16'h23d9, 16'h23d4, 16'h23cf, 16'h23ca, 16'h23c5, 16'h23c0, 16'h23bb, 16'h23b6, 16'h23b1, 16'h23ac, 16'h23a7, 16'h23a2, 16'h239d, 16'h2398, 16'h2393, 16'h238e, 16'h2389, 16'h2384, 16'h237f, 16'h237a, 16'h2375, 16'h2370, 16'h236b, 16'h2366, 16'h2361, 16'h235c, 16'h2357, 16'h2352, 16'h234d, 16'h2348, 16'h2343, 16'h233e, 16'h2339, 16'h2334, 16'h232f, 16'h232a, 16'h2325, 16'h2320, 16'h231b, 16'h2316, 16'h2311, 16'h230c, 16'h2307, 16'h2302, 16'h22fd},
                                 {16'h22f8, 16'h22f3, 16'h22ee, 16'h22e9, 16'h22e4, 16'h22df, 16'h22da, 16'h22d5, 16'h22d0, 16'h22cb, 16'h22c6, 16'h22c1, 16'h22bc, 16'h22b7, 16'h22b2, 16'h22ad, 16'h22a8, 16'h22a3, 16'h229e, 16'h2299, 16'h2294, 16'h228f, 16'h228a, 16'h2285, 16'h2280, 16'h227b, 16'h2276, 16'h2271, 16'h226c, 16'h2267, 16'h2262, 16'h225d, 16'h2258, 16'h2253, 16'h224e, 16'h2249, 16'h2244, 16'h223f, 16'h223a, 16'h2235, 16'h2230, 16'h222b, 16'h2226, 16'h2221, 16'h221c, 16'h2217, 16'h2212, 16'h220d, 16'h2208, 16'h2203, 16'h21fe, 16'h21f9, 16'h21f4, 16'h21ef, 16'h21ea, 16'h21e5, 16'h21e0, 16'h21db, 16'h21d6, 16'h21d1, 16'h21cc, 16'h21c7, 16'h21c2, 16'h21bd},
                                 {16'h21b8, 16'h21b3, 16'h21ae, 16'h21a9, 16'h21a4, 16'h219f, 16'h219a, 16'h2195, 16'h2190, 16'h218b, 16'h2186, 16'h2181, 16'h217c, 16'h2177, 16'h2172, 16'h216d, 16'h2168, 16'h2163, 16'h215e, 16'h2159, 16'h2154, 16'h214f, 16'h214a, 16'h2145, 16'h2140, 16'h213b, 16'h2136, 16'h2131, 16'h212c, 16'h2127, 16'h2122, 16'h211d, 16'h2118, 16'h2113, 16'h210e, 16'h2109, 16'h2104, 16'h20ff, 16'h20fa, 16'h20f5, 16'h20f0, 16'h20eb, 16'h20e6, 16'h20e1, 16'h20dc, 16'h20d7, 16'h20d2, 16'h20cd, 16'h20c8, 16'h20c3, 16'h20be, 16'h20b9, 16'h20b4, 16'h20af, 16'h20aa, 16'h20a5, 16'h20a0, 16'h209b, 16'h2096, 16'h2091, 16'h208c, 16'h2087, 16'h2082, 16'h207d},
                                 {16'h2078, 16'h2073, 16'h206e, 16'h2069, 16'h2064, 16'h205f, 16'h205a, 16'h2055, 16'h2050, 16'h204b, 16'h2046, 16'h2041, 16'h203c, 16'h2037, 16'h2032, 16'h202d, 16'h2028, 16'h2023, 16'h201e, 16'h2019, 16'h2014, 16'h200f, 16'h200a, 16'h2005, 16'h2000, 16'h1ffb, 16'h1ff6, 16'h1ff1, 16'h1fec, 16'h1fe7, 16'h1fe2, 16'h1fdd, 16'h1fd8, 16'h1fd3, 16'h1fce, 16'h1fc9, 16'h1fc4, 16'h1fbf, 16'h1fba, 16'h1fb5, 16'h1fb0, 16'h1fab, 16'h1fa6, 16'h1fa1, 16'h1f9c, 16'h1f97, 16'h1f92, 16'h1f8d, 16'h1f88, 16'h1f83, 16'h1f7e, 16'h1f79, 16'h1f74, 16'h1f6f, 16'h1f6a, 16'h1f65, 16'h1f60, 16'h1f5b, 16'h1f56, 16'h1f51, 16'h1f4c, 16'h1f47, 16'h1f42, 16'h1f3d},
                                 {16'h1f38, 16'h1f33, 16'h1f2e, 16'h1f29, 16'h1f24, 16'h1f1f, 16'h1f1a, 16'h1f15, 16'h1f10, 16'h1f0b, 16'h1f06, 16'h1f01, 16'h1efc, 16'h1ef7, 16'h1ef2, 16'h1eed, 16'h1ee8, 16'h1ee3, 16'h1ede, 16'h1ed9, 16'h1ed4, 16'h1ecf, 16'h1eca, 16'h1ec5, 16'h1ec0, 16'h1ebb, 16'h1eb6, 16'h1eb1, 16'h1eac, 16'h1ea7, 16'h1ea2, 16'h1e9d, 16'h1e98, 16'h1e93, 16'h1e8e, 16'h1e89, 16'h1e84, 16'h1e7f, 16'h1e7a, 16'h1e75, 16'h1e70, 16'h1e6b, 16'h1e66, 16'h1e61, 16'h1e5c, 16'h1e57, 16'h1e52, 16'h1e4d, 16'h1e48, 16'h1e43, 16'h1e3e, 16'h1e39, 16'h1e34, 16'h1e2f, 16'h1e2a, 16'h1e25, 16'h1e20, 16'h1e1b, 16'h1e16, 16'h1e11, 16'h1e0c, 16'h1e07, 16'h1e02, 16'h1dfd},
                                 {16'h1df8, 16'h1df4, 16'h1df0, 16'h1dec, 16'h1de8, 16'h1de4, 16'h1de0, 16'h1ddc, 16'h1dd8, 16'h1dd4, 16'h1dd0, 16'h1dcc, 16'h1dc8, 16'h1dc4, 16'h1dc0, 16'h1dbc, 16'h1db8, 16'h1db4, 16'h1db0, 16'h1dac, 16'h1da8, 16'h1da4, 16'h1da0, 16'h1d9c, 16'h1d98, 16'h1d94, 16'h1d90, 16'h1d8c, 16'h1d88, 16'h1d84, 16'h1d80, 16'h1d7c, 16'h1d78, 16'h1d74, 16'h1d70, 16'h1d6c, 16'h1d68, 16'h1d64, 16'h1d60, 16'h1d5c, 16'h1d58, 16'h1d54, 16'h1d50, 16'h1d4c, 16'h1d48, 16'h1d44, 16'h1d40, 16'h1d3c, 16'h1d38, 16'h1d34, 16'h1d30, 16'h1d2c, 16'h1d28, 16'h1d24, 16'h1d20, 16'h1d1c, 16'h1d18, 16'h1d14, 16'h1d10, 16'h1d0c, 16'h1d08, 16'h1d04, 16'h1d00, 16'h1cfc},
                                 {16'h1cf8, 16'h1cf4, 16'h1cf0, 16'h1cec, 16'h1ce8, 16'h1ce4, 16'h1ce0, 16'h1cdc, 16'h1cd8, 16'h1cd4, 16'h1cd0, 16'h1ccc, 16'h1cc8, 16'h1cc4, 16'h1cc0, 16'h1cbc, 16'h1cb8, 16'h1cb4, 16'h1cb0, 16'h1cac, 16'h1ca8, 16'h1ca4, 16'h1ca0, 16'h1c9c, 16'h1c98, 16'h1c94, 16'h1c90, 16'h1c8c, 16'h1c88, 16'h1c84, 16'h1c80, 16'h1c7c, 16'h1c78, 16'h1c74, 16'h1c70, 16'h1c6c, 16'h1c68, 16'h1c64, 16'h1c60, 16'h1c5c, 16'h1c58, 16'h1c54, 16'h1c50, 16'h1c4c, 16'h1c48, 16'h1c44, 16'h1c40, 16'h1c3c, 16'h1c38, 16'h1c34, 16'h1c30, 16'h1c2c, 16'h1c28, 16'h1c24, 16'h1c20, 16'h1c1c, 16'h1c18, 16'h1c14, 16'h1c10, 16'h1c0c, 16'h1c08, 16'h1c04, 16'h1c00, 16'h1bfc},
                                 {16'h1bf8, 16'h1bf4, 16'h1bf0, 16'h1bec, 16'h1be8, 16'h1be4, 16'h1be0, 16'h1bdc, 16'h1bd8, 16'h1bd4, 16'h1bd0, 16'h1bcc, 16'h1bc8, 16'h1bc4, 16'h1bc0, 16'h1bbc, 16'h1bb8, 16'h1bb4, 16'h1bb0, 16'h1bac, 16'h1ba8, 16'h1ba4, 16'h1ba0, 16'h1b9c, 16'h1b98, 16'h1b94, 16'h1b90, 16'h1b8c, 16'h1b88, 16'h1b84, 16'h1b80, 16'h1b7c, 16'h1b78, 16'h1b74, 16'h1b70, 16'h1b6c, 16'h1b68, 16'h1b64, 16'h1b60, 16'h1b5c, 16'h1b58, 16'h1b54, 16'h1b50, 16'h1b4c, 16'h1b48, 16'h1b44, 16'h1b40, 16'h1b3c, 16'h1b38, 16'h1b34, 16'h1b30, 16'h1b2c, 16'h1b28, 16'h1b24, 16'h1b20, 16'h1b1c, 16'h1b18, 16'h1b14, 16'h1b10, 16'h1b0c, 16'h1b08, 16'h1b04, 16'h1b00, 16'h1afc},
                                 {16'h1af8, 16'h1af4, 16'h1af0, 16'h1aec, 16'h1ae8, 16'h1ae4, 16'h1ae0, 16'h1adc, 16'h1ad8, 16'h1ad4, 16'h1ad0, 16'h1acc, 16'h1ac8, 16'h1ac4, 16'h1ac0, 16'h1abc, 16'h1ab8, 16'h1ab4, 16'h1ab0, 16'h1aac, 16'h1aa8, 16'h1aa4, 16'h1aa0, 16'h1a9c, 16'h1a98, 16'h1a94, 16'h1a90, 16'h1a8c, 16'h1a88, 16'h1a84, 16'h1a80, 16'h1a7c, 16'h1a78, 16'h1a74, 16'h1a70, 16'h1a6c, 16'h1a68, 16'h1a64, 16'h1a60, 16'h1a5c, 16'h1a58, 16'h1a54, 16'h1a50, 16'h1a4c, 16'h1a48, 16'h1a44, 16'h1a40, 16'h1a3c, 16'h1a38, 16'h1a34, 16'h1a30, 16'h1a2c, 16'h1a28, 16'h1a24, 16'h1a20, 16'h1a1c, 16'h1a18, 16'h1a14, 16'h1a10, 16'h1a0c, 16'h1a08, 16'h1a04, 16'h1a00, 16'h19fc},
                                 {16'h19f8, 16'h19f4, 16'h19f0, 16'h19ec, 16'h19e8, 16'h19e4, 16'h19e0, 16'h19dc, 16'h19d8, 16'h19d4, 16'h19d0, 16'h19cc, 16'h19c8, 16'h19c4, 16'h19c0, 16'h19bc, 16'h19b8, 16'h19b4, 16'h19b0, 16'h19ac, 16'h19a8, 16'h19a4, 16'h19a0, 16'h199c, 16'h1998, 16'h1994, 16'h1990, 16'h198c, 16'h1988, 16'h1984, 16'h1980, 16'h197c, 16'h1978, 16'h1974, 16'h1970, 16'h196c, 16'h1968, 16'h1964, 16'h1960, 16'h195c, 16'h1958, 16'h1954, 16'h1950, 16'h194c, 16'h1948, 16'h1944, 16'h1940, 16'h193c, 16'h1938, 16'h1934, 16'h1930, 16'h192c, 16'h1928, 16'h1924, 16'h1920, 16'h191c, 16'h1918, 16'h1914, 16'h1910, 16'h190c, 16'h1908, 16'h1904, 16'h1900, 16'h18fc},
                                 {16'h18f8, 16'h18f4, 16'h18f0, 16'h18ec, 16'h18e8, 16'h18e4, 16'h18e0, 16'h18dc, 16'h18d8, 16'h18d4, 16'h18d0, 16'h18cc, 16'h18c8, 16'h18c4, 16'h18c0, 16'h18bc, 16'h18b8, 16'h18b4, 16'h18b0, 16'h18ac, 16'h18a8, 16'h18a4, 16'h187f, 16'h1872, 16'h1865, 16'h1858, 16'h184b, 16'h183e, 16'h1831, 16'h1824, 16'h1817, 16'h180a, 16'h17fd, 16'h17f0, 16'h17e3, 16'h17d6, 16'h17c9, 16'h17bc, 16'h17af, 16'h17a2, 16'h1795, 16'h1788, 16'h177b, 16'h176e, 16'h1761, 16'h1754, 16'h1747, 16'h173a, 16'h172d, 16'h1720, 16'h1713, 16'h1706, 16'h16f9, 16'h16ec, 16'h16df, 16'h16d2, 16'h16c5, 16'h16b8, 16'h16ab, 16'h169e, 16'h1691, 16'h1684, 16'h1677, 16'h166a},
                                 {16'h165d, 16'h1650, 16'h1643, 16'h1636, 16'h1629, 16'h161c, 16'h160f, 16'h1602, 16'h15f5, 16'h15e8, 16'h15db, 16'h15ce, 16'h15c1, 16'h15b4, 16'h15a7, 16'h159a, 16'h158d, 16'h1580, 16'h1573, 16'h1566, 16'h1559, 16'h154c, 16'h153f, 16'h1532, 16'h1525, 16'h1518, 16'h150b, 16'h14fe, 16'h14f1, 16'h14e4, 16'h14d7, 16'h14ca, 16'h14bd, 16'h14b0, 16'h14a3, 16'h1496, 16'h1489, 16'h147c, 16'h146f, 16'h1462, 16'h1455, 16'h1448, 16'h143b, 16'h142e, 16'h1421, 16'h1414, 16'h1407, 16'h13fa, 16'h13ed, 16'h13e0, 16'h13d3, 16'h13c6, 16'h13b9, 16'h13ac, 16'h139f, 16'h1392, 16'h1385, 16'h1378, 16'h136b, 16'h135e, 16'h1351, 16'h1344, 16'h1337, 16'h132a},
                                 {16'h131d, 16'h1310, 16'h1303, 16'h12f6, 16'h12e9, 16'h12dc, 16'h12cf, 16'h12c2, 16'h12b5, 16'h12a8, 16'h129b, 16'h128e, 16'h1281, 16'h1274, 16'h1267, 16'h125a, 16'h124d, 16'h1240, 16'h1233, 16'h1226, 16'h1219, 16'h120c, 16'h11ff, 16'h11f2, 16'h11e5, 16'h11d8, 16'h11cb, 16'h11be, 16'h11b1, 16'h11a4, 16'h1197, 16'h118a, 16'h117d, 16'h1170, 16'h1163, 16'h1156, 16'h1149, 16'h113c, 16'h112f, 16'h1122, 16'h1115, 16'h1108, 16'h10fb, 16'h10ee, 16'h10e1, 16'h10d4, 16'h10c7, 16'h10ba, 16'h10ad, 16'h10a0, 16'h1093, 16'h1086, 16'h1079, 16'h106c, 16'h105f, 16'h1052, 16'h1045, 16'h1038, 16'h102b, 16'h101e, 16'h1011, 16'h1004, 16'h0ff7, 16'h0fea},
                                 {16'h0fdd, 16'h0fd0, 16'h0fc3, 16'h0fb6, 16'h0fa9, 16'h0f9c, 16'h0f8f, 16'h0f82, 16'h0f75, 16'h0f68, 16'h0f5b, 16'h0f4e, 16'h0f41, 16'h0f34, 16'h0f27, 16'h0f1a, 16'h0f0d, 16'h0f00, 16'h0ef3, 16'h0ee6, 16'h0ed9, 16'h0ecc, 16'h0ebf, 16'h0eb2, 16'h0ea5, 16'h0e98, 16'h0e8b, 16'h0e7e, 16'h0e71, 16'h0e64, 16'h0e57, 16'h0e4a, 16'h0e3d, 16'h0e30, 16'h0e23, 16'h0e16, 16'h0e09, 16'h0dfc, 16'h0def, 16'h0de2, 16'h0dd5, 16'h0dc8, 16'h0dbb, 16'h0dae, 16'h0da1, 16'h0d94, 16'h0d87, 16'h0d7a, 16'h0d6d, 16'h0d60, 16'h0d53, 16'h0d46, 16'h0d39, 16'h0d2c, 16'h0d1f, 16'h0d12, 16'h0d05, 16'h0cf8, 16'h0ceb, 16'h0cde, 16'h0cd1, 16'h0cc4, 16'h0cb7, 16'h0caa},
                                 {16'h0c9d, 16'h0c90, 16'h0c83, 16'h0c76, 16'h0c69, 16'h0c5c, 16'h0c4f, 16'h0c42, 16'h0c35, 16'h0c28, 16'h0c1b, 16'h0c0e, 16'h0c01, 16'h0bf4, 16'h0be7, 16'h0bda, 16'h0bcd, 16'h0bc0, 16'h0bb3, 16'h0ba6, 16'h0b99, 16'h0b8c, 16'h0b7f, 16'h0b72, 16'h0b65, 16'h0b58, 16'h0b4b, 16'h0b3e, 16'h0b31, 16'h0b24, 16'h0b17, 16'h0b0a, 16'h0afd, 16'h0af0, 16'h0ae3, 16'h0ad6, 16'h0ac9, 16'h0abc, 16'h1a87, 16'h19b9, 16'h19ad, 16'h19a1, 16'h1995, 16'h1989, 16'h197d, 16'h1971, 16'h1965, 16'h1959, 16'h194d, 16'h1941, 16'h1935, 16'h1929, 16'h191d, 16'h1911, 16'h1905, 16'h18f9, 16'h18ed, 16'h18e1, 16'h18d5, 16'h18c9, 16'h18bd, 16'h18b1, 16'h18a5, 16'h1899},
                                 {16'h188d, 16'h1881, 16'h1875, 16'h1869, 16'h185d, 16'h1851, 16'h1845, 16'h1839, 16'h182d, 16'h1821, 16'h1815, 16'h1809, 16'h17fd, 16'h17f1, 16'h17e5, 16'h17d9, 16'h17cd, 16'h17c1, 16'h17b5, 16'h17a9, 16'h179d, 16'h1791, 16'h1785, 16'h1779, 16'h176d, 16'h1761, 16'h1755, 16'h1749, 16'h173d, 16'h1731, 16'h1725, 16'h1719, 16'h170d, 16'h1701, 16'h16f5, 16'h16e9, 16'h16dd, 16'h16d1, 16'h16c5, 16'h16b9, 16'h16ad, 16'h16a1, 16'h1695, 16'h1689, 16'h167d, 16'h1671, 16'h1665, 16'h1659, 16'h164d, 16'h1641, 16'h1635, 16'h1629, 16'h161d, 16'h1611, 16'h1605, 16'h15f9, 16'h15ed, 16'h15e1, 16'h15d5, 16'h15c9, 16'h15bd, 16'h15b1, 16'h15a5, 16'h1599},
                                 {16'h158d, 16'h1581, 16'h1575, 16'h1569, 16'h155d, 16'h1551, 16'h1545, 16'h1539, 16'h152d, 16'h1521, 16'h1515, 16'h1509, 16'h14fd, 16'h14f1, 16'h14e5, 16'h14d9, 16'h14cd, 16'h14c1, 16'h14b5, 16'h14a9, 16'h149d, 16'h1491, 16'h1485, 16'h1479, 16'h146d, 16'h1461, 16'h1455, 16'h1449, 16'h143d, 16'h1431, 16'h1425, 16'h1419, 16'h140d, 16'h1401, 16'h13f5, 16'h13e9, 16'h13dd, 16'h13d1, 16'h13c5, 16'h13b9, 16'h13ad, 16'h13a1, 16'h1395, 16'h1389, 16'h137d, 16'h1371, 16'h1365, 16'h1359, 16'h134d, 16'h1341, 16'h1335, 16'h1329, 16'h131d, 16'h1311, 16'h1305, 16'h12f9, 16'h12ed, 16'h12e1, 16'h12d5, 16'h12c9, 16'h12bd, 16'h12b1, 16'h12a5, 16'h1299},
                                 {16'h128d, 16'h1281, 16'h1275, 16'h1269, 16'h125d, 16'h1251, 16'h1245, 16'h1239, 16'h122d, 16'h1221, 16'h1215, 16'h1209, 16'h11fd, 16'h11f1, 16'h11e5, 16'h11d9, 16'h11cd, 16'h11c1, 16'h11b5, 16'h11a9, 16'h119d, 16'h1191, 16'h1185, 16'h1179, 16'h116d, 16'h1161, 16'h1155, 16'h1149, 16'h113d, 16'h1131, 16'h1125, 16'h1119, 16'h110d, 16'h1101, 16'h10f5, 16'h10e9, 16'h10dd, 16'h10d1, 16'h10c5, 16'h10b9, 16'h10ad, 16'h10a1, 16'h1095, 16'h1089, 16'h107d, 16'h1071, 16'h1065, 16'h1059, 16'h104d, 16'h1041, 16'h1035, 16'h1029, 16'h101d, 16'h1011, 16'h1005, 16'h0ff9, 16'h0fed, 16'h0fe1, 16'h0fd5, 16'h0fc9, 16'h0fbd, 16'h0fb1, 16'h0fa5, 16'h0f99},
                                 {16'h0f8d, 16'h0f81, 16'h0f75, 16'h0f69, 16'h0f5d, 16'h0f51, 16'h0f45, 16'h0f39, 16'h0f2d, 16'h0f21, 16'h0f15, 16'h0f09, 16'h0efd, 16'h0ef1, 16'h0ee5, 16'h0ed9, 16'h0ecd, 16'h0ec1, 16'h0eb5, 16'h0ea9, 16'h0e9d, 16'h0e91, 16'h0e85, 16'h0e79, 16'h0e6d, 16'h0e61, 16'h0e55, 16'h0e49, 16'h0e3d, 16'h0e31, 16'h0e25, 16'h0e19, 16'h0e0d, 16'h0e01, 16'h0df5, 16'h0de9, 16'h0ddd, 16'h0dd1, 16'h0dc5, 16'h0db9, 16'h0dad, 16'h0da1, 16'h0d95, 16'h0d89, 16'h0d7d, 16'h0d71, 16'h0d65, 16'h0d59, 16'h0d4d, 16'h0d41, 16'h0d35, 16'h0d29, 16'h0d1d, 16'h0d11, 16'h0d05, 16'h0cf9, 16'h0ced, 16'h0ce1, 16'h0cd5, 16'h0cc9, 16'h0cbd, 16'h0cb1, 16'h0ca5, 16'h0c99},
                                 {16'h0c8d, 16'h0c81, 16'h0c75, 16'h0c69, 16'h0c5d, 16'h0c51, 16'h0c45, 16'h0c39, 16'h0c2d, 16'h0c21, 16'h0c15, 16'h0c09, 16'h0bfd, 16'h0bf1, 16'h0be5, 16'h0bd9, 16'h0bcd, 16'h0bc1, 16'h0bb5, 16'h0ba9, 16'h0b9d, 16'h0b91, 16'h0b85, 16'h0b79, 16'h0b6d, 16'h0b61, 16'h0b55, 16'h0b49, 16'h0b3d, 16'h0b31, 16'h0b25, 16'h0b19, 16'h0b0d, 16'h0b01, 16'h0af5, 16'h0ae9, 16'h0add, 16'h0ad1, 16'h0ac5, 16'h0ab9, 16'h0aad, 16'h0aa1, 16'h0a95, 16'h0a89, 16'h0a7d, 16'h0a71, 16'h0a65, 16'h0a59, 16'h0a4d, 16'h0a41, 16'h0a35, 16'h0a29, 16'h0a1d, 16'h0a11, 16'h0a05, 16'h09f9, 16'h09ed, 16'h09e1, 16'h09d5, 16'h09c9, 16'h09bd, 16'h09b1, 16'h09a5, 16'h0999},
                                 {16'h098d, 16'h0981, 16'h0975, 16'h0969, 16'h095d, 16'h0951, 16'h0945, 16'h0939, 16'h092d, 16'h0921, 16'h0915, 16'h0909, 16'h08fd, 16'h08f1, 16'h08e5, 16'h08d9, 16'h08cd, 16'h08c1, 16'h08b5, 16'h08a9, 16'h089d, 16'h0891, 16'h0885, 16'h0879, 16'h086d, 16'h0861, 16'h0855, 16'h0849, 16'h083d, 16'h0831, 16'h0825, 16'h0819, 16'h080d, 16'h0801, 16'h07f5, 16'h07e9, 16'h07dd, 16'h07d1, 16'h07c5, 16'h07b9, 16'h07ad, 16'h07a1, 16'h0795, 16'h081d, 16'h08a9, 16'h0935, 16'h09c1, 16'h0a4d, 16'h0ad9, 16'h0b65, 16'h0bf1, 16'h0c7d, 16'h0d09, 16'h0d95, 16'h0e21, 16'h0ead, 16'h0f39, 16'h0fc5, 16'h1051, 16'h10dd, 16'h1169, 16'h11f5, 16'h1281, 16'h130d},
                                 {16'h1399, 16'h1425, 16'h14b1, 16'h153d, 16'h15c9, 16'h1655, 16'h16e1, 16'h176d, 16'h17f9, 16'h1885, 16'h1911, 16'h199d, 16'h1a29, 16'h1ab5, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41},
                                 {16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41},
                                 {16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41},
                                 {16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41},
                                 {16'h1b41, 16'h1b41, 16'h1b41, 16'h1b41, 16'h1b40, 16'h1b3f, 16'h1b3e, 16'h1b3d, 16'h1b3c, 16'h1b3b, 16'h1b3a, 16'h1b39, 16'h1b38, 16'h1b37, 16'h1b36, 16'h1b35, 16'h1b34, 16'h1b33, 16'h1b32, 16'h1b31, 16'h1b30, 16'h1b2f, 16'h1b2e, 16'h1b2d, 16'h1b2c, 16'h1b2b, 16'h1b2a, 16'h1b29, 16'h1b28, 16'h1b27, 16'h1b26, 16'h1b25, 16'h1b24, 16'h1b23, 16'h1b22, 16'h1b21, 16'h1b20, 16'h1b1f, 16'h1b1e, 16'h1b1d, 16'h1b1c, 16'h1b1b, 16'h1b1a, 16'h1b19, 16'h1b18, 16'h1b17, 16'h1b16, 16'h1b15, 16'h1b14, 16'h1b13, 16'h1b12, 16'h1b11, 16'h1b10, 16'h1b0f, 16'h1b0e, 16'h1b0d, 16'h1b0c, 16'h1b0b, 16'h1b0a, 16'h1b09, 16'h1b08, 16'h1b07, 16'h1b06, 16'h1b05},
                                 {16'h1ac7, 16'h1ab7, 16'h1aa7, 16'h1a97, 16'h1a87, 16'h1a77, 16'h1a67, 16'h1a57, 16'h1a47, 16'h1a37, 16'h1a27, 16'h1a17, 16'h1a07, 16'h19f7, 16'h19e7, 16'h19d7, 16'h19c7, 16'h19b7, 16'h19a7, 16'h1997, 16'h1987, 16'h1977, 16'h1967, 16'h1957, 16'h1947, 16'h1937, 16'h1927, 16'h1917, 16'h1907, 16'h18f7, 16'h18e7, 16'h18d7, 16'h18c7, 16'h18b7, 16'h18a7, 16'h1897, 16'h1887, 16'h1877, 16'h1867, 16'h1857, 16'h1847, 16'h1837, 16'h1827, 16'h1817, 16'h1807, 16'h17f7, 16'h17e7, 16'h17d7, 16'h17c7, 16'h17b7, 16'h17a7, 16'h1797, 16'h1787, 16'h1777, 16'h1767, 16'h1757, 16'h1747, 16'h1737, 16'h1727, 16'h1717, 16'h1707, 16'h16f7, 16'h16e7, 16'h16d7},
                                 {16'h16c7, 16'h16b7, 16'h16a7, 16'h1697, 16'h1687, 16'h1677, 16'h1667, 16'h1657, 16'h1647, 16'h1637, 16'h1627, 16'h1617, 16'h1607, 16'h15f7, 16'h15e7, 16'h15d7, 16'h15c7, 16'h15b7, 16'h15a7, 16'h1597, 16'h1587, 16'h1577, 16'h1567, 16'h1557, 16'h1547, 16'h1537, 16'h1527, 16'h1517, 16'h1507, 16'h14f7, 16'h14e7, 16'h14d7, 16'h14c7, 16'h14b7, 16'h14a7, 16'h1497, 16'h1487, 16'h1477, 16'h1467, 16'h1457, 16'h1447, 16'h1437, 16'h1427, 16'h1417, 16'h1407, 16'h13f7, 16'h13e7, 16'h13d7, 16'h13c7, 16'h13b7, 16'h13a7, 16'h1397, 16'h1387, 16'h1377, 16'h1367, 16'h1357, 16'h1347, 16'h1337, 16'h1327, 16'h1317, 16'h1307, 16'h12f7, 16'h12e7, 16'h12d7},
                                 {16'h12c7, 16'h12b7, 16'h12a7, 16'h1297, 16'h1287, 16'h1277, 16'h1267, 16'h1257, 16'h1247, 16'h1237, 16'h1227, 16'h1217, 16'h1207, 16'h11f7, 16'h11e7, 16'h11d7, 16'h11c7, 16'h11b7, 16'h11a7, 16'h1197, 16'h1187, 16'h1177, 16'h1167, 16'h1157, 16'h1147, 16'h1137, 16'h1127, 16'h1117, 16'h1107, 16'h10f7, 16'h10e7, 16'h10d7, 16'h10c7, 16'h10b7, 16'h10a7, 16'h1097, 16'h1087, 16'h1077, 16'h1067, 16'h1057, 16'h1047, 16'h1037, 16'h1027, 16'h1017, 16'h1007, 16'h0ff7, 16'h0fe7, 16'h0fd7, 16'h0fc7, 16'h0fb7, 16'h0fa7, 16'h0f97, 16'h0f87, 16'h0f77, 16'h0f67, 16'h0f57, 16'h0f47, 16'h0f37, 16'h0f27, 16'h0f17, 16'h0f07, 16'h0ef7, 16'h0ee7, 16'h0ed7},
                                 {16'h0ec7, 16'h0eb7, 16'h0ea7, 16'h0e97, 16'h0e87, 16'h0e77, 16'h0e67, 16'h0e57, 16'h0e47, 16'h0e37, 16'h0e27, 16'h0e17, 16'h0e07, 16'h0df7, 16'h0de7, 16'h0dd7, 16'h0dc7, 16'h0db7, 16'h0da7, 16'h0d97, 16'h0d87, 16'h0d77, 16'h0d67, 16'h0d57, 16'h0d47, 16'h0d37, 16'h0d27, 16'h0d17, 16'h0d07, 16'h0cf7, 16'h0ce7, 16'h0cd7, 16'h0cc7, 16'h0cb7, 16'h0ca7, 16'h0c97, 16'h0c87, 16'h0c77, 16'h0c67, 16'h0c57, 16'h0c47, 16'h0c37, 16'h0c27, 16'h0c17, 16'h0c07, 16'h0bf7, 16'h0be7, 16'h0bd7, 16'h0bc7, 16'h0bb7, 16'h0ba7, 16'h0b97, 16'h0b87, 16'h0b77, 16'h0b67, 16'h0b57, 16'h0b47, 16'h0b37, 16'h0b27, 16'h0b17, 16'h0b07, 16'h0af7, 16'h0ae7, 16'h0ad7},
                                 {16'h0ac7, 16'h0ab7, 16'h0aa7, 16'h0a97, 16'h0a87, 16'h0a77, 16'h0a77, 16'h0a77, 16'h0a8e, 16'h0ab9, 16'h0ae4, 16'h0b0f, 16'h0b3a, 16'h0b65, 16'h0b90, 16'h0bbb, 16'h0be6, 16'h0c11, 16'h0c3c, 16'h0c67, 16'h0c92, 16'h0cbd, 16'h0ce8, 16'h0d13, 16'h0d3e, 16'h0d69, 16'h0d94, 16'h0dbf, 16'h0dea, 16'h0e15, 16'h0e40, 16'h0e6b, 16'h0e96, 16'h0ec1, 16'h0eec, 16'h0f17, 16'h0f42, 16'h0f6d, 16'h0f98, 16'h0fc3, 16'h0fee, 16'h1019, 16'h1044, 16'h106f, 16'h109a, 16'h10c5, 16'h10f0, 16'h111b, 16'h1146, 16'h1171, 16'h119c, 16'h11c7, 16'h11f2, 16'h121d, 16'h1248, 16'h1273, 16'h129e, 16'h12c9, 16'h12f4, 16'h131f, 16'h134a, 16'h1375, 16'h13a0, 16'h13cb},
                                 {16'h13f6, 16'h1421, 16'h144c, 16'h1477, 16'h14a2, 16'h14cd, 16'h14f8, 16'h1523, 16'h154e, 16'h1579, 16'h15a4, 16'h15cf, 16'h15fa, 16'h1625, 16'h1650, 16'h167b, 16'h16a6, 16'h16d1, 16'h16fc, 16'h1727, 16'h1752, 16'h177d, 16'h17a8, 16'h17d3, 16'h17fe, 16'h1829, 16'h1854, 16'h187f, 16'h18aa, 16'h18d5, 16'h1900, 16'h192b, 16'h1956, 16'h1981, 16'h19ac, 16'h19d7, 16'h1a02, 16'h1a2d, 16'h1a58, 16'h1a83, 16'h1aae, 16'h1ad9, 16'h1b04, 16'h1b2f, 16'h1b5a, 16'h1b85, 16'h1bb0, 16'h1bdb, 16'h1c06, 16'h1c31, 16'h1c5c, 16'h1c87, 16'h1cb2, 16'h1cdd, 16'h1d08, 16'h1d33, 16'h1d5e, 16'h1d89, 16'h1db4, 16'h1ddf, 16'h1e0a, 16'h1e35, 16'h1e60, 16'h1e8b},
                                 {16'h1eb6, 16'h1ee1, 16'h1f0c, 16'h1f37, 16'h1f62, 16'h1f8d, 16'h1fb8, 16'h1fe3, 16'h200e, 16'h2039, 16'h2064, 16'h208f, 16'h20ba, 16'h20e5, 16'h2110, 16'h213b, 16'h2166, 16'h2191, 16'h21bc, 16'h21e7, 16'h2212, 16'h223d, 16'h2268, 16'h2293, 16'h22be, 16'h22e9, 16'h2314, 16'h233f, 16'h236a, 16'h2395, 16'h23c0, 16'h23eb, 16'h2416, 16'h2441, 16'h246c, 16'h2497, 16'h24c2, 16'h24ed, 16'h2518, 16'h2543, 16'h256e, 16'h2599, 16'h25c4, 16'h25ef, 16'h261a, 16'h2645, 16'h2670, 16'h269b, 16'h26c6, 16'h26f1, 16'h271c, 16'h2747, 16'h2772, 16'h279d, 16'h27c8, 16'h27f3, 16'h281e, 16'h2849, 16'h2874, 16'h289f, 16'h28ca, 16'h28f5, 16'h2920, 16'h294b},
                                 {16'h2976, 16'h29a1, 16'h29cc, 16'h29f7, 16'h2a22, 16'h2a4d, 16'h2a78, 16'h2aa3, 16'h2ace, 16'h2af9, 16'h2b24, 16'h2b4f, 16'h2b7a, 16'h2ba5, 16'h2bd0, 16'h2bfb, 16'h2c26, 16'h2c51, 16'h2c7c, 16'h2ca7, 16'h2cd2, 16'h2cfd, 16'h2d28, 16'h2d53, 16'h2d7e, 16'h2da9, 16'h2dd4, 16'h2dff, 16'h2e2a, 16'h2e55, 16'h2e80, 16'h2eab, 16'h2ed6, 16'h2f01, 16'h2f2c, 16'h2f57, 16'h2f82, 16'h2fad, 16'h2fd8, 16'h3003, 16'h302e, 16'h3059, 16'h3084, 16'h30af, 16'h30da, 16'h3105, 16'h3130, 16'h315b, 16'h3186, 16'h31b1, 16'h31dc, 16'h3207, 16'h3232, 16'h325d, 16'h3288, 16'h32b3, 16'h32de, 16'h3309, 16'h3334, 16'h335f, 16'h338a, 16'h33b5, 16'h33e0, 16'h340b},
                                 {16'h3436, 16'h3461, 16'h348c, 16'h34b7, 16'h34e2, 16'h350d, 16'h3538, 16'h3563, 16'h358e, 16'h35b9, 16'h35e4, 16'h360f, 16'h363a, 16'h3665, 16'h3690, 16'h36bb, 16'h36e6, 16'h3711, 16'h373c, 16'h3767, 16'h3792, 16'h37bd, 16'h37e8, 16'h3813, 16'h383e, 16'h3869, 16'h3894, 16'h38bf, 16'h38ea, 16'h3915, 16'h3940, 16'h396b, 16'h3996, 16'h39c1, 16'h39ec, 16'h3a17, 16'h3a42, 16'h3a6d, 16'h3a98, 16'h3ac3, 16'h3aee, 16'h3b19, 16'h3b44, 16'h3b6f, 16'h3b9a, 16'h3bc5, 16'h3bf0, 16'h3c1b, 16'h3c46, 16'h3c71, 16'h3c9c, 16'h3cc7, 16'h3cf2, 16'h3d1d, 16'h3d48, 16'h3d73, 16'h3d9e, 16'h3dc9, 16'h3df4, 16'h3e1f, 16'h3e50, 16'h3e50, 16'h3e20, 16'h3de9},
                                 {16'h3db2, 16'h3d7b, 16'h3d44, 16'h3d0d, 16'h3cd6, 16'h3c9f, 16'h3c68, 16'h3c31, 16'h3bfa, 16'h3bc3, 16'h3b8c, 16'h3b55, 16'h3b1e, 16'h3ae7, 16'h3ab0, 16'h3a79, 16'h3a42, 16'h3a0b, 16'h39d4, 16'h399d, 16'h3966, 16'h392f, 16'h38f8, 16'h38c1, 16'h388a, 16'h3853, 16'h381c, 16'h37e5, 16'h37ae, 16'h3777, 16'h3740, 16'h3709, 16'h36d2, 16'h369b, 16'h3664, 16'h362d, 16'h35f6, 16'h35bf, 16'h3588, 16'h3551, 16'h351a, 16'h34e3, 16'h34ac, 16'h3475, 16'h343e, 16'h3407, 16'h33d0, 16'h3399, 16'h3362, 16'h332b, 16'h32f4, 16'h32bd, 16'h3286, 16'h324f, 16'h3218, 16'h31e1, 16'h31aa, 16'h3173, 16'h313c, 16'h3105, 16'h30ce, 16'h3097, 16'h3060, 16'h3029},
                                 {16'h2ff2, 16'h2fbb, 16'h2f84, 16'h2f4d, 16'h2f16, 16'h2edf, 16'h2ea8, 16'h2e71, 16'h2e3a, 16'h2e03, 16'h2dcc, 16'h2d95, 16'h2d5e, 16'h2d27, 16'h2cf0, 16'h2cb9, 16'h2c82, 16'h2c4b, 16'h2c14, 16'h2bdd, 16'h2ba6, 16'h2b6f, 16'h2b38, 16'h2b01, 16'h2aca, 16'h2a93, 16'h2a5c, 16'h2a25, 16'h29ee, 16'h29b7, 16'h2980, 16'h2949, 16'h2912, 16'h28db, 16'h28a4, 16'h286d, 16'h2836, 16'h27ff, 16'h27c8, 16'h2791, 16'h275a, 16'h2723, 16'h26ec, 16'h26b5, 16'h267e, 16'h2647, 16'h2610, 16'h25d9, 16'h25a2, 16'h256b, 16'h2534, 16'h24fd, 16'h24c6, 16'h248f, 16'h2458, 16'h2421, 16'h23ea, 16'h23b3, 16'h237c, 16'h2345, 16'h230e, 16'h22d7, 16'h22a0, 16'h2269},
                                 {16'h2232, 16'h21fb, 16'h21c4, 16'h218d, 16'h2156, 16'h211f, 16'h20e8, 16'h20b1, 16'h207a, 16'h2043, 16'h200c, 16'h1fd5, 16'h1f9e, 16'h1f67, 16'h1f30, 16'h1ef9, 16'h1ec2, 16'h1e8b, 16'h1e54, 16'h1e1d, 16'h1de6, 16'h1daf, 16'h1d78, 16'h1d41, 16'h1d0a, 16'h1cd3, 16'h1c9c, 16'h1c65, 16'h1c2e, 16'h1bf7, 16'h1bc0, 16'h1b89, 16'h1b52, 16'h1b1b, 16'h1ae4, 16'h1aad, 16'h1a76, 16'h1a3f, 16'h1a08, 16'h19d1, 16'h199a, 16'h1963, 16'h192c, 16'h18f5, 16'h18be, 16'h1887, 16'h1850, 16'h1819, 16'h17e2, 16'h17ab, 16'h1774, 16'h173d, 16'h1706, 16'h16cf, 16'h1698, 16'h1661, 16'h162a, 16'h15f3, 16'h15bc, 16'h1585, 16'h154e, 16'h1517, 16'h14e0, 16'h14a9},
                                 {16'h1472, 16'h143b, 16'h1404, 16'h13cd, 16'h13cd, 16'h13cd, 16'h13cd, 16'h13cd, 16'h13cd, 16'h13cd, 16'h13cd, 16'h13cd, 16'h13cd, 16'h13cd, 16'h13cd, 16'h13cd, 16'h13cd, 16'h13cd, 16'h13cd, 16'h13cd, 16'h13cd, 16'h13cd, 16'h13cd, 16'h13cd, 16'h13da, 16'h13e7, 16'h13f4, 16'h1401, 16'h140e, 16'h141b, 16'h1428, 16'h1435, 16'h1442, 16'h144f, 16'h145c, 16'h1469, 16'h1476, 16'h1483, 16'h1490, 16'h149d, 16'h14aa, 16'h14b7, 16'h14c4, 16'h14d1, 16'h14de, 16'h14eb, 16'h14f8, 16'h1505, 16'h1512, 16'h151f, 16'h152c, 16'h1539, 16'h1546, 16'h1553, 16'h1560, 16'h156d, 16'h157a, 16'h1587, 16'h1594, 16'h15a1, 16'h15ae, 16'h15bb, 16'h15c8, 16'h15d5},
                                 {16'h15e2, 16'h15ef, 16'h15fc, 16'h1609, 16'h1616, 16'h1623, 16'h1630, 16'h163d, 16'h164a, 16'h1657, 16'h1664, 16'h1671, 16'h167e, 16'h168b, 16'h1698, 16'h16a5, 16'h16b2, 16'h16bf, 16'h16cc, 16'h16d9, 16'h16e6, 16'h16f3, 16'h1700, 16'h170d, 16'h171a, 16'h1727, 16'h1734, 16'h1741, 16'h174e, 16'h175b, 16'h1768, 16'h1775, 16'h1782, 16'h178f, 16'h179c, 16'h17a9, 16'h17b6, 16'h17c3, 16'h17d0, 16'h17dd, 16'h17ea, 16'h17f7, 16'h1804, 16'h1811, 16'h181e, 16'h182b, 16'h1838, 16'h1845, 16'h1852, 16'h185f, 16'h186c, 16'h1879, 16'h1886, 16'h1893, 16'h18a0, 16'h18ad, 16'h18ba, 16'h18c7, 16'h18d4, 16'h18e1, 16'h18ee, 16'h18fb, 16'h1908, 16'h1915},
                                 {16'h1922, 16'h192f, 16'h193c, 16'h1949, 16'h1956, 16'h1963, 16'h1970, 16'h197d, 16'h198a, 16'h1997, 16'h19a4, 16'h19b1, 16'h19be, 16'h19cb, 16'h19d8, 16'h19e5, 16'h19f2, 16'h19ff, 16'h1a0c, 16'h1a19, 16'h1a26, 16'h1a33, 16'h1a40, 16'h1a4d, 16'h1a5a, 16'h1a67, 16'h1a74, 16'h1a81, 16'h1a8e, 16'h1a9b, 16'h1aa8, 16'h1ab5, 16'h1ac2, 16'h1acf, 16'h1adc, 16'h1ae9, 16'h1af6, 16'h1b03, 16'h1b10, 16'h1b1d, 16'h1b2a, 16'h1b37, 16'h1b44, 16'h1b51, 16'h1b5e, 16'h1b6b, 16'h1b78, 16'h1b85, 16'h1b92, 16'h1b9f, 16'h1bac, 16'h1bb9, 16'h1bc6, 16'h1bd3, 16'h1be0, 16'h1bed, 16'h1bfa, 16'h1c07, 16'h1c14, 16'h1c21, 16'h1c2e, 16'h1c3b, 16'h1c48, 16'h1c55},
                                 {16'h1c62, 16'h1c6f, 16'h1c7c, 16'h1c89, 16'h1c96, 16'h1ca3, 16'h1cb0, 16'h1cbd, 16'h1cca, 16'h1cd7, 16'h1ce4, 16'h1cf1, 16'h1cfe, 16'h1d0b, 16'h1d18, 16'h1d25, 16'h1d32, 16'h1d3f, 16'h1d4c, 16'h1d59, 16'h1d66, 16'h1d73, 16'h1d80, 16'h1d8d, 16'h1d9a, 16'h1da7, 16'h1db4, 16'h1dc1, 16'h1dce, 16'h1ddb, 16'h1de8, 16'h1df5, 16'h1e02, 16'h1e0f, 16'h1e1c, 16'h1e29, 16'h1e36, 16'h1e43, 16'h1e50, 16'h1e5d, 16'h1e6a, 16'h1e77, 16'h1e84, 16'h1e91, 16'h1e9e, 16'h1eab, 16'h1eb8, 16'h1ec5, 16'h1ed2, 16'h1edf, 16'h1eec, 16'h1ef9, 16'h1f06, 16'h1f13, 16'h1f20, 16'h1f2d, 16'h1f3a, 16'h1f47, 16'h1f54, 16'h1f61, 16'h1f6e, 16'h1f7b, 16'h1f88, 16'h1f95},
                                 {16'h1fa2, 16'h1faf, 16'h1fbc, 16'h1fc9, 16'h1fd6, 16'h1fe3, 16'h1ff0, 16'h1ffd, 16'h200a, 16'h2017, 16'h2024, 16'h2031, 16'h203e, 16'h204b, 16'h2058, 16'h2065, 16'h2072, 16'h207f, 16'h208c, 16'h2099, 16'h20a6, 16'h20b3, 16'h20c0, 16'h20cd, 16'h20da, 16'h20e7, 16'h20f4, 16'h2101, 16'h210e, 16'h211b, 16'h2128, 16'h2135, 16'h2142, 16'h214f, 16'h215c, 16'h2169, 16'h2176, 16'h2183, 16'h2190, 16'h219d, 16'h21aa, 16'h21b7, 16'h21c4, 16'h21d1, 16'h21de, 16'h21eb, 16'h21f8, 16'h2205, 16'h2212, 16'h221f, 16'h222c, 16'h2239, 16'h2246, 16'h2253, 16'h2260, 16'h226d, 16'h227a, 16'h2287, 16'h2294, 16'h22a1, 16'h22ae, 16'h22bb, 16'h22c8, 16'h22d5},
                                 {16'h22e2, 16'h22ef, 16'h22fc, 16'h2309, 16'h2316, 16'h2323, 16'h2330, 16'h233d, 16'h234a, 16'h2357, 16'h2364, 16'h2371, 16'h237e, 16'h238b, 16'h2398, 16'h23a5, 16'h23b2, 16'h23bf, 16'h23cc, 16'h23d9, 16'h23e6, 16'h23f3, 16'h2400, 16'h240d, 16'h241a, 16'h2427, 16'h2434, 16'h2441, 16'h244e, 16'h245b, 16'h2468, 16'h2475, 16'h2482, 16'h248f, 16'h249c, 16'h24a9, 16'h24b6, 16'h24c3, 16'h24d0, 16'h24dd, 16'h24ea, 16'h24f7, 16'h2504, 16'h2511, 16'h251e, 16'h252b, 16'h2538, 16'h2545, 16'h2552, 16'h255f, 16'h256c, 16'h2579, 16'h2586, 16'h2593, 16'h25a0, 16'h25ad, 16'h25ba, 16'h25c7, 16'h25d4, 16'h25e1, 16'h25ee, 16'h25fb, 16'h2608, 16'h2615},
                                 {16'h2622, 16'h262f, 16'h263c, 16'h2649, 16'h2656, 16'h2663, 16'h2670, 16'h267d, 16'h268a, 16'h2697, 16'h26a4, 16'h26b1, 16'h26be, 16'h26cb, 16'h26d8, 16'h26e5, 16'h26f2, 16'h26ff, 16'h270c, 16'h2719, 16'h2726, 16'h2733, 16'h2740, 16'h274d, 16'h275a, 16'h2767, 16'h2774, 16'h2781, 16'h278e, 16'h279b, 16'h27a8, 16'h27b5, 16'h27c2, 16'h27cf, 16'h27dc, 16'h27e9, 16'h27f6, 16'h2803, 16'h2810, 16'h281d, 16'h282a, 16'h2837, 16'h2844, 16'h2851, 16'h285e, 16'h286b, 16'h2878, 16'h2885, 16'h2892, 16'h289f, 16'h28ac, 16'h28b9, 16'h28c6, 16'h28d3, 16'h28e0, 16'h28ed, 16'h28fa, 16'h2907, 16'h2914, 16'h2921, 16'h292e, 16'h293b, 16'h2948, 16'h2955},
                                 {16'h2962, 16'h296f, 16'h297c, 16'h2989, 16'h2996, 16'h29a3, 16'h29b0, 16'h29bd, 16'h29ca, 16'h29d7, 16'h29e4, 16'h29f1, 16'h29fe, 16'h2a0b, 16'h2a18, 16'h2a25, 16'h2a32, 16'h2a3f, 16'h2a4c, 16'h2a59, 16'h2a66, 16'h2a73, 16'h2a80, 16'h2a8d, 16'h2a9a, 16'h2aa7, 16'h2ab4, 16'h2ac1, 16'h2ace, 16'h2adb, 16'h2ae8, 16'h2af5, 16'h2b02, 16'h2b0f, 16'h2b1c, 16'h2b29, 16'h2b36, 16'h2b43, 16'h2b50, 16'h2b5d, 16'h2b6a, 16'h2b77, 16'h2b84, 16'h2b91, 16'h2b9e, 16'h2bab, 16'h2bb8, 16'h2bc5, 16'h2bd2, 16'h2bdf, 16'h2bec, 16'h2bf9, 16'h2c06, 16'h2c13, 16'h2c20, 16'h2c2d, 16'h2c3a, 16'h2c47, 16'h2c54, 16'h2c61, 16'h2c6e, 16'h2c7b, 16'h2c88, 16'h2c95},
                                 {16'h2ca2, 16'h2caf, 16'h2cbc, 16'h2cc9, 16'h2cd6, 16'h2ce3, 16'h2cf0, 16'h2cfd, 16'h2d0a, 16'h2d17, 16'h2d24, 16'h2d31, 16'h2d3e, 16'h2d4b, 16'h2d58, 16'h2d65, 16'h2d72, 16'h2d7f, 16'h2d8c, 16'h2d99, 16'h2da6, 16'h2db3, 16'h2dc0, 16'h2dcd, 16'h2dda, 16'h2de7, 16'h2df4, 16'h2e01, 16'h2e0e, 16'h2e1b, 16'h2e28, 16'h2e35, 16'h2e42, 16'h2e4f, 16'h2e5c, 16'h2e69, 16'h2e76, 16'h2e83, 16'h2e90, 16'h2e9d, 16'h2eaa, 16'h2eb7, 16'h2ec4, 16'h2ed1, 16'h2ede, 16'h2eeb, 16'h2ef8, 16'h2f05, 16'h2f12, 16'h2f1f, 16'h2f2c, 16'h2f39, 16'h2f46, 16'h2f53, 16'h2f60, 16'h2f6d, 16'h2f7a, 16'h2f87, 16'h2f94, 16'h2fa1, 16'h2fae, 16'h2fbb, 16'h2fc8, 16'h2fd5},
                                 {16'h2fe2, 16'h2fef, 16'h2ffc, 16'h3009, 16'h3016, 16'h3023, 16'h3030, 16'h303d, 16'h304a, 16'h3057, 16'h3064, 16'h3071, 16'h307e, 16'h308b, 16'h3098, 16'h30a5, 16'h30b2, 16'h30bf, 16'h30cc, 16'h30d9, 16'h30e6, 16'h30f3, 16'h3100, 16'h310d, 16'h311a, 16'h3127, 16'h3134, 16'h3141, 16'h314e, 16'h315b, 16'h3168, 16'h3175, 16'h3182, 16'h318f, 16'h319c, 16'h31a9, 16'h2056, 16'h20da, 16'h20ee, 16'h2102, 16'h2116, 16'h212a, 16'h213e, 16'h2152, 16'h2166, 16'h217a, 16'h218e, 16'h21a2, 16'h21b6, 16'h21ca, 16'h21de, 16'h21f2, 16'h2206, 16'h221a, 16'h222e, 16'h2242, 16'h2256, 16'h226a, 16'h227e, 16'h2292, 16'h22a6, 16'h22ba, 16'h22ce, 16'h22e2},
                                 {16'h22f6, 16'h230a, 16'h231e, 16'h2332, 16'h2346, 16'h235a, 16'h236e, 16'h2382, 16'h2396, 16'h23aa, 16'h23be, 16'h23d2, 16'h23e6, 16'h23fa, 16'h240e, 16'h2422, 16'h2436, 16'h244a, 16'h245e, 16'h2472, 16'h2486, 16'h249a, 16'h24ae, 16'h24c2, 16'h24d6, 16'h24ea, 16'h24fe, 16'h2512, 16'h2526, 16'h253a, 16'h254e, 16'h2562, 16'h2576, 16'h258a, 16'h259e, 16'h25b2, 16'h25c6, 16'h25da, 16'h25ee, 16'h2602, 16'h2616, 16'h262a, 16'h263e, 16'h2652, 16'h2666, 16'h267a, 16'h268e, 16'h26a2, 16'h26b6, 16'h26ca, 16'h26de, 16'h26f2, 16'h2706, 16'h271a, 16'h272e, 16'h2742, 16'h2756, 16'h276a, 16'h277e, 16'h2792, 16'h27a6, 16'h27ba, 16'h27ce, 16'h27e2},
                                 {16'h27f6, 16'h280a, 16'h281e, 16'h2832, 16'h2846, 16'h285a, 16'h286e, 16'h2882, 16'h2896, 16'h28aa, 16'h28be, 16'h28d2, 16'h28e6, 16'h28fa, 16'h290e, 16'h2922, 16'h2936, 16'h294a, 16'h295e, 16'h2972, 16'h2986, 16'h299a, 16'h29ae, 16'h29c2, 16'h29d6, 16'h29ea, 16'h29fe, 16'h2a12, 16'h2a26, 16'h2a3a, 16'h2a4e, 16'h2a62, 16'h2a76, 16'h2a8a, 16'h2a9e, 16'h2ab2, 16'h2ac6, 16'h2ada, 16'h2aee, 16'h2b02, 16'h2b16, 16'h2b2a, 16'h2b3e, 16'h2b52, 16'h2b66, 16'h2b7a, 16'h2b8e, 16'h2ba2, 16'h2bb6, 16'h2bca, 16'h2bde, 16'h2bf2, 16'h2c06, 16'h2c1a, 16'h2c2e, 16'h2c42, 16'h2c56, 16'h2c6a, 16'h2c7e, 16'h2c92, 16'h2ca6, 16'h2cba, 16'h2cce, 16'h2ce2},
                                 {16'h2cf6, 16'h2d0a, 16'h2d1e, 16'h2d32, 16'h2d46, 16'h2d5a, 16'h2d6e, 16'h2d82, 16'h2d96, 16'h2daa, 16'h2dbe, 16'h2dd2, 16'h2de6, 16'h2dfa, 16'h2e0e, 16'h2e22, 16'h2e36, 16'h2e4a, 16'h2e5e, 16'h2e72, 16'h2e86, 16'h2e9a, 16'h2eae, 16'h2ec2, 16'h2ed6, 16'h2eea, 16'h2efe, 16'h2f12, 16'h2f26, 16'h2f3a, 16'h2f4e, 16'h2f62, 16'h2f76, 16'h2f8a, 16'h2f9e, 16'h2fb2, 16'h2fc6, 16'h2fda, 16'h2fee, 16'h3002, 16'h3016, 16'h302a, 16'h303e, 16'h3052, 16'h3066, 16'h307a, 16'h308e, 16'h30a2, 16'h30b6, 16'h30ca, 16'h30de, 16'h30f2, 16'h3106, 16'h311a, 16'h312e, 16'h3142, 16'h3156, 16'h316a, 16'h317e, 16'h3192, 16'h31a6, 16'h31ba, 16'h31ce, 16'h31e2},
                                 {16'h31f6, 16'h320a, 16'h321e, 16'h3232, 16'h3246, 16'h325a, 16'h326e, 16'h3282, 16'h3296, 16'h32aa, 16'h32be, 16'h32d2, 16'h32e6, 16'h32fa, 16'h330e, 16'h3322, 16'h3336, 16'h334a, 16'h335e, 16'h3372, 16'h3386, 16'h339a, 16'h33ae, 16'h33c2, 16'h33d6, 16'h33ea, 16'h33fe, 16'h3412, 16'h3426, 16'h343a, 16'h344e, 16'h3462, 16'h3476, 16'h348a, 16'h349e, 16'h34b2, 16'h34c6, 16'h34da, 16'h34ee, 16'h3502, 16'h3516, 16'h352a, 16'h353e, 16'h3552, 16'h3566, 16'h357a, 16'h358e, 16'h35a2, 16'h35b6, 16'h35ca, 16'h35de, 16'h35f2, 16'h3606, 16'h361a, 16'h362e, 16'h3642, 16'h3656, 16'h366a, 16'h367e, 16'h3692, 16'h36a6, 16'h36ba, 16'h36ce, 16'h36e2},
                                 {16'h36f6, 16'h370a, 16'h371e, 16'h3732, 16'h3746, 16'h375a, 16'h376e, 16'h3782, 16'h3796, 16'h37aa, 16'h37be, 16'h37d2, 16'h37e6, 16'h37fa, 16'h380e, 16'h3822, 16'h3836, 16'h384a, 16'h385e, 16'h3872, 16'h3886, 16'h389a, 16'h38ae, 16'h38c2, 16'h38c2, 16'h38c2, 16'h38c2, 16'h38c2, 16'h38bb, 16'h389a, 16'h3879, 16'h3858, 16'h3837, 16'h3816, 16'h37f5, 16'h37d4, 16'h37b3, 16'h3792, 16'h3771, 16'h3750, 16'h372f, 16'h370e, 16'h36ed, 16'h36cc, 16'h36ab, 16'h368a, 16'h3669, 16'h3648, 16'h3627, 16'h3606, 16'h35e5, 16'h35c4, 16'h35a3, 16'h3582, 16'h3561, 16'h3540, 16'h351f, 16'h34fe, 16'h34dd, 16'h34bc, 16'h349b, 16'h347a, 16'h3459, 16'h3438},
                                 {16'h3417, 16'h33f6, 16'h33d5, 16'h33b4, 16'h3393, 16'h3372, 16'h3351, 16'h3330, 16'h330f, 16'h32ee, 16'h32cd, 16'h32ac, 16'h328b, 16'h326a, 16'h3249, 16'h3228, 16'h3207, 16'h31e6, 16'h31c5, 16'h31a4, 16'h3183, 16'h3162, 16'h3141, 16'h3120, 16'h30ff, 16'h30de, 16'h30bd, 16'h309c, 16'h307b, 16'h305a, 16'h3039, 16'h3018, 16'h2ff7, 16'h2fd6, 16'h2fb5, 16'h2f94, 16'h2f73, 16'h2f52, 16'h2f31, 16'h2f10, 16'h2eef, 16'h2ece, 16'h2ead, 16'h2e8c, 16'h2e6b, 16'h2e4a, 16'h2e29, 16'h2e08, 16'h2de7, 16'h2dc6, 16'h2da5, 16'h2d84, 16'h2d63, 16'h2d42, 16'h2d21, 16'h2d00, 16'h2cdf, 16'h2cbe, 16'h2c9d, 16'h2c7c, 16'h2c5b, 16'h2c3a, 16'h2c19, 16'h2bf8},
                                 {16'h2bd7, 16'h2bb6, 16'h2b95, 16'h2b74, 16'h2b53, 16'h2b32, 16'h2b11, 16'h2af0, 16'h2acf, 16'h2aae, 16'h2a8d, 16'h2a6c, 16'h2a4b, 16'h2a2a, 16'h2a09, 16'h29e8, 16'h29c7, 16'h29a6, 16'h2985, 16'h2964, 16'h2943, 16'h2922, 16'h2901, 16'h28e0, 16'h28bf, 16'h289e, 16'h287d, 16'h285c, 16'h283b, 16'h281a, 16'h27f9, 16'h27d8, 16'h27b7, 16'h2796, 16'h2775, 16'h2754, 16'h2733, 16'h2712, 16'h26f1, 16'h26d0, 16'h26af, 16'h268e, 16'h266d, 16'h264c, 16'h262b, 16'h260a, 16'h25e9, 16'h25c8, 16'h25a7, 16'h2586, 16'h2565, 16'h2544, 16'h2523, 16'h2502, 16'h24e1, 16'h24c0, 16'h249f, 16'h247e, 16'h245d, 16'h243c, 16'h241b, 16'h23fa, 16'h23d9, 16'h23b8},
                                 {16'h2397, 16'h2376, 16'h2355, 16'h2334, 16'h2313, 16'h22f2, 16'h22d1, 16'h22b0, 16'h228f, 16'h226e, 16'h224d, 16'h222c, 16'h220b, 16'h21ea, 16'h21c9, 16'h21a8, 16'h2187, 16'h2166, 16'h2145, 16'h2124, 16'h2103, 16'h20e2, 16'h20c1, 16'h20a0, 16'h207f, 16'h205e, 16'h203d, 16'h201c, 16'h1ffb, 16'h1fda, 16'h1fb9, 16'h1f98, 16'h1f77, 16'h1f56, 16'h1f35, 16'h1f14, 16'h1ef3, 16'h1ed2, 16'h1eb1, 16'h1e90, 16'h1e6f, 16'h1e4e, 16'h1e2d, 16'h1e0c, 16'h1deb, 16'h1dca, 16'h1da9, 16'h1d88, 16'h1d67, 16'h1d46, 16'h1d25, 16'h1d04, 16'h1ce3, 16'h1cc2, 16'h1ca1, 16'h1c80, 16'h1c5f, 16'h1c3e, 16'h1c1d, 16'h1bfc, 16'h1bdb, 16'h1bba, 16'h1b99, 16'h1b78},
                                 {16'h1b57, 16'h1b36, 16'h1b15, 16'h1af4, 16'h1ad3, 16'h1ab2, 16'h1a91, 16'h1a70, 16'h1a4f, 16'h1a2e, 16'h1a0d, 16'h19ec, 16'h19cb, 16'h19aa, 16'h1989, 16'h1968, 16'h1947, 16'h1926, 16'h1905, 16'h18e4, 16'h18c3, 16'h18a2, 16'h1881, 16'h1860, 16'h183f, 16'h181e, 16'h17fd, 16'h17dc, 16'h17bb, 16'h179a, 16'h1779, 16'h1758, 16'h1737, 16'h1716, 16'h16f5, 16'h16d4, 16'h16b3, 16'h1692, 16'h1671, 16'h1650, 16'h162f, 16'h160e, 16'h15ed, 16'h15cc, 16'h15ab, 16'h158a, 16'h1569, 16'h1548, 16'h1527, 16'h1506, 16'h14e5, 16'h14c4, 16'h14a3, 16'h1482, 16'h1461, 16'h1440, 16'h141f, 16'h13fe, 16'h13dd, 16'h13bc, 16'h139b, 16'h137a, 16'h1359, 16'h1338},
                                 {16'h1317, 16'h12f6, 16'h12d5, 16'h12b4, 16'h1293, 16'h1272, 16'h1251, 16'h1230, 16'h120f, 16'h11ee, 16'h11cd, 16'h11ac, 16'h118b, 16'h116a, 16'h1149, 16'h1128, 16'h1107, 16'h10e6, 16'h10c5, 16'h10a4, 16'h1083, 16'h1062, 16'h1041, 16'h1020, 16'h0fff, 16'h0fde, 16'h0fbd, 16'h0f9c, 16'h0f7b, 16'h0f5a, 16'h0f39, 16'h0f18, 16'h0ef7, 16'h0ed6, 16'h0eb5, 16'h0e94, 16'h0401, 16'h0401, 16'h0401, 16'h0401, 16'h0401, 16'h0401, 16'h03ff, 16'h03fc, 16'h03f9, 16'h03f6, 16'h03f3, 16'h03f0, 16'h03ed, 16'h03ea, 16'h03e7, 16'h03e4, 16'h03e1, 16'h03de, 16'h03db, 16'h03d8, 16'h03d5, 16'h03d2, 16'h03cf, 16'h03cc, 16'h03c9, 16'h03c6, 16'h03c3, 16'h03c0},
                                 {16'h03bd, 16'h03ba, 16'h03b7, 16'h03b4, 16'h03b1, 16'h03ae, 16'h03ab, 16'h03a8, 16'h03a5, 16'h03a2, 16'h039f, 16'h039c, 16'h0399, 16'h0396, 16'h0393, 16'h0390, 16'h038d, 16'h038a, 16'h0387, 16'h0384, 16'h0381, 16'h037e, 16'h037b, 16'h0378, 16'h0375, 16'h0372, 16'h036f, 16'h036c, 16'h0369, 16'h0366, 16'h0363, 16'h0360, 16'h035d, 16'h035a, 16'h0357, 16'h0354, 16'h0351, 16'h034e, 16'h034b, 16'h0348, 16'h0345, 16'h0342, 16'h033f, 16'h033c, 16'h0339, 16'h0336, 16'h0333, 16'h0330, 16'h032d, 16'h032a, 16'h0327, 16'h0324, 16'h0321, 16'h031e, 16'h031b, 16'h0318, 16'h0315, 16'h0312, 16'h030f, 16'h030c, 16'h0309, 16'h0306, 16'h0303, 16'h0300},
                                 {16'h02fd, 16'h02fa, 16'h02f7, 16'h02f4, 16'h02f1, 16'h02ee, 16'h02eb, 16'h02e8, 16'h02e5, 16'h02e2, 16'h02df, 16'h02dc, 16'h02d9, 16'h02d6, 16'h02d3, 16'h02d0, 16'h02cd, 16'h02ca, 16'h02c7, 16'h02c4, 16'h02c1, 16'h02be, 16'h02bb, 16'h02b8, 16'h02b5, 16'h02b2, 16'h02af, 16'h02ac, 16'h02a9, 16'h02a6, 16'h02a3, 16'h02a0, 16'h029d, 16'h029a, 16'h0297, 16'h0294, 16'h0291, 16'h028e, 16'h028b, 16'h0288, 16'h0285, 16'h0282, 16'h027f, 16'h027c, 16'h0279, 16'h0276, 16'h0273, 16'h0270, 16'h026d, 16'h026a, 16'h0267, 16'h0264, 16'h0261, 16'h025e, 16'h025b, 16'h0258, 16'h0255, 16'h0252, 16'h024f, 16'h024c, 16'h0249, 16'h0246, 16'h0243, 16'h0240},
                                 {16'h023d, 16'h023a, 16'h0237, 16'h0234, 16'h0231, 16'h022e, 16'h022b, 16'h0228, 16'h0225, 16'h0222, 16'h021f, 16'h021c, 16'h0219, 16'h0216, 16'h0213, 16'h0210, 16'h020d, 16'h020a, 16'h0207, 16'h0204, 16'h0201, 16'h01fe, 16'h01fb, 16'h01f8, 16'h01f5, 16'h01f2, 16'h01ef, 16'h01ec, 16'h01e9, 16'h01e6, 16'h01e3, 16'h01e0, 16'h01dd, 16'h01da, 16'h01d7, 16'h01d4, 16'h01d1, 16'h01ce, 16'h01cb, 16'h01c8, 16'h01c5, 16'h01c2, 16'h01bf, 16'h01bc, 16'h01b9, 16'h01b6, 16'h01b3, 16'h01b0, 16'h01ad, 16'h01aa, 16'h01a7, 16'h01a4, 16'h01a1, 16'h019e, 16'h019b, 16'h0198, 16'h0195, 16'h0192, 16'h018f, 16'h018c, 16'h0189, 16'h0186, 16'h0183, 16'h0180},
                                 {16'h017d, 16'h017a, 16'h0177, 16'h0174, 16'h0171, 16'h016e, 16'h016b, 16'h0168, 16'h0165, 16'h0162, 16'h015f, 16'h015c, 16'h0159, 16'h0156, 16'h0153, 16'h0150, 16'h014d, 16'h014a, 16'h0147, 16'h0144, 16'h0141, 16'h013e, 16'h013b, 16'h0138, 16'h0135, 16'h0132, 16'h012f, 16'h012c, 16'h0129, 16'h0126, 16'h0123, 16'h0120, 16'h011d, 16'h011a, 16'h0117, 16'h0114, 16'h0111, 16'h010e, 16'h010b, 16'h0108, 16'h0105, 16'h0102, 16'h00ff, 16'h00fc, 16'h00f9, 16'h00f6, 16'h00f3, 16'h00f0, 16'h00ed, 16'h00ea, 16'h00e7, 16'h00e4, 16'h00e1, 16'h00de, 16'h00db, 16'h00d8, 16'h00d5, 16'h00d2, 16'h00cf, 16'h00cc, 16'h00c9, 16'h00c6, 16'h00c3, 16'h00c0},
                                 {16'h00bd, 16'h00ba, 16'h00b7, 16'h00b4, 16'h00b1, 16'h00ae, 16'h00ab, 16'h00a8, 16'h00a5, 16'h00a2, 16'h009f, 16'h009c, 16'h0099, 16'h0096, 16'h0093, 16'h0090, 16'h008d, 16'h008a, 16'h0087, 16'h0084, 16'h0081, 16'h007e, 16'h007b, 16'h0078, 16'h0075, 16'h0072, 16'h006f, 16'h006c, 16'h0069, 16'h0066, 16'h0063, 16'h0060, 16'h005d, 16'h005a, 16'h0057, 16'h0054, 16'h0051, 16'h004e, 16'h004b, 16'h0048, 16'h0045, 16'h0042, 16'h003f, 16'h003c, 16'h0039, 16'h0036, 16'h0033, 16'h0030, 16'h002d, 16'h002a, 16'h0027, 16'h0024, 16'h0021, 16'h001e, 16'h001b, 16'h0018, 16'h0015, 16'h0012, 16'h000f, 16'h000c, 16'h0009, 16'h0006, 16'h0003, 16'h0000}};
    /*
    FOLLOWING PATH: (time,val,slope)
    (0, 0, 3) --> (347, 1025, 2707) --> (348, 3732, 33) --> (680, 14530, -20) --> (987, 8278, 4435) --> (988, 12713, -13)
    (1596, 5069, 55) --> (1795, 15952, -49) --> (1796, 15903, -43) --> (2106, 2679, 16) --> (2368, 6917, 1)
    (2673, 6977, -140) --> (2709, 1941, 12) --> (3097, 6791, -4043) --> (3098, 2748, 13) --> (3370, 6308, 4)
    (3712, 7677, 5) --> (4039, 9221, -59) --> (4186, 492, 8) --> (4466, 2610, 7440) --> (4467, 10050, -23)
    (4716, 4305, -23) --> (4830, 1645, 1) --> (5069, 1680, 17) --> (5662, 11647, -8) --> (5917, 9619, -57)
    (5957, 7324, 24) --> (6276, 14974, -3) --> (6668, 13631, 6) --> (6827, 14599, -3) --> (6931, 14245, -14)
    (7203, 10468, 19) --> (7426, 14647, -39) --> (7754, 1979, 8765) --> (7755, 10744, -28) --> (8039, 2704, 1)
    (8250, 2925, 16) --> (8658, 9337, -177) --> (8707, 679, 24) --> (9078, 9762, -52) --> (9094, 8928, 15)
    (9249, 11185, 6) --> (9783, 14268, -620) --> (9784, 13648, -28) --> (10141, 3803, 17) --> (10382, 7807, 53)
    (10425, 10075, 10) --> (10966, 15594, -60) --> (11171, 3241, 34) --> (11371, 10084, -8432) --> (11372, 1652, 45)
    (11515, 8023, -8) --> (12070, 3804, 2) --> (12316, 4387, -4) --> (12562, 3429, 3587) --> (12563, 7016, -19)
    (12877, 1036, 6) --> (12913, 1267, 26) --> (13379, 13418, -33) --> (13559, 7427, 22) --> (13936, 15737, -9)
    (14027, 14910, -103) --> (14166, 624, 1) --> (14598, 1044, 36) --> (14872, 10893, -1) --> (15144, 10869, -31)
    (15412, 2431, 0)
    */
    top_level tl(.clk(clk),
                 .sys_rst(rst),
                 .dac0_rdy(dac0_rdy),
                 .dac_batch(dac_batch),
                 .valid_dac_batch(valid_dac_batch),
                 .pl_rstn(pl_rstn),
                 .raddr_packet(raddr_packet),
                 .raddr_valid_packet(raddr_valid_packet),
                 .waddr_packet(waddr_packet),
                 .waddr_valid_packet(waddr_valid_packet),
                 .wdata_packet(wdata_packet),
                 .wdata_valid_packet(wdata_valid_packet),
                 .ps_wresp_rdy(ps_wresp_rdy),
                 .ps_read_rdy(ps_read_rdy),
                 .wresp_out(wresp_out),
                 .rresp_out(rresp_out),
                 .wresp_valid_out(wresp_valid_out),
                 .rresp_valid_out(rresp_valid_out),
                 .rdata_packet(rdata_packet),
                 .rdata_valid_out(rdata_valid_out),
                 .pwl_tdata(pwl_tdata),
                 .pwl_tkeep(pwl_tkeep),
                 .pwl_tlast(pwl_tlast),
                 .pwl_tvalid(pwl_tvalid),
                 .pwl_tready(pwl_tready));

    oscillate_sig #(.DELAY (10))
    dac_rdy_oscillator(.clk(clk), .rst(rst), .long_on(1'b0),
                       .osc_sig_out(dac0_rdy));
    oscillate_sig #(.DELAY (25))
    read_rdy_oscillator(.clk(clk), .rst(rst), .long_on(1'b0),
                        .osc_sig_out(ps_read_rdy));
    oscillate_sig #(.DELAY (30))
    wresp_rdy_oscillator(.clk(clk), .rst(rst), .long_on(1'b0),
                        .osc_sig_out(ps_wresp_rdy));
    generate
        for (genvar i = 0; i < `BATCH_SAMPLES; i++) begin: batch_splices
            data_splicer #(.DATA_WIDTH(`BATCH_WIDTH), .SPLICE_WIDTH(`SAMPLE_WIDTH))
            dac_out_splice(.data(dac_batch),
                           .i(int'(i)),
                           .spliced_data(dac_samples[i]));
        end
    endgenerate

    assign curr_expected_batch = expected_batches[exp_i];
    assign checked_full_wave = (pwlTestState == VERIFY) && (valid_dac_batch) && (exp_i == (tl.sys.dac_intf.pwl_gen.wave_lines_stored-1)); 
    assign curr_expected_batch = expected_batches[exp_i];
    always_comb begin
        if (test_num == 0) 
            test_check = {tl.sys.rst,tl.sys.rst};
        else if (test_num == 1)
            test_check = (rdata_valid_out && ps_read_rdy && testState == TEST)? {rdata_packet == `MAX_ILA_BURST_SIZE,1'b1} : 0; 
        else if (test_num == 2) begin
            if (valid_dac_batch) begin
                for (int i = 0; i < `BATCH_WIDTH; i++) error_vec[i] = dac_samples[i] != curr_expected_batch[i]; 
            end else error_vec = 0; 
            test_check = (valid_dac_batch)? {dac_batch == curr_expected_batch,1'b1} : 0; 
        end
        else {test_check, error_vec} = 0; 
    end

    always_ff @(posedge clk) begin
        if (rst || panic) begin
            if (panic) begin
                testState <= DONE;
                kill_tb <= 1; 
                panic <= 0;
            end else begin
                testState <= IDLE;
                {testsPassed,testsFailed, kill_tb} <= 0; 
                {done, timer} <= 0;
                test_num <= STARTING_TEST; 

                {raddr_packet, waddr_packet, wdata_packet} <= 0;
                {raddr_valid_packet, waddr_valid_packet, wdata_valid_packet} <= 0; 
                {pwl_tlast, pwl_tdata, pwl_tvalid} <= 0;
                {dma_i,exp_i,send_dma_buff,run_pwl,periods} <= 0;
                pwlTestState <= IDLE_PWL; 
            end
        end else begin
            case(pwlTestState)
                IDLE_PWL: begin 
                    if (send_dma_buff) begin
                        pwl_tvalid <= 1; 
                        pwl_tdata = dma_buff[0];
                        pwl_tlast <= 0; 
                        dma_i <= 1; 
                        pwlTestState <= SEND_BUFF; 
                    end
                    if (run_pwl) begin
                        {pwl_tlast, pwl_tdata, pwl_tvalid,dma_i} <= 0;
                        {exp_i, periods} <= 0;
                        pwlTestState <= VERIFY;  
                    end
                end  
                SEND_BUFF: begin
                    if (dma_i < BUFF_LEN) begin
                        if (pwl_tready) begin
                            pwl_tdata = dma_buff[dma_i];
                            if (dma_i == BUFF_LEN-1) pwl_tlast <= 1; 
                            dma_i <= dma_i + 1;
                        end 
                    end
                    else if (dma_i == BUFF_LEN && pwl_tready) begin
                        {pwl_tlast, pwl_tdata, pwl_tvalid} <= 0;
                        dma_i <= 0;
                        pwlTestState <= VERIFY;  
                    end
                end 
                VERIFY: begin
                    if (periods == PERIODS_TO_CHECK) begin
                        {exp_i, periods} <= 0;
                        pwlTestState <= IDLE_PWL;
                    end else if (checked_full_wave) begin
                        periods <= periods + 1;
                        exp_i <= 0; 
                    end else if (valid_dac_batch) exp_i <= exp_i + 1; 
                end 
            endcase

            case(testState)
                IDLE: begin 
                    if (start) testState <= TEST; 
                    if (done) done <= 0; 
                end 
                TEST: begin
                    // Write to reset
                    if (test_num == 0) begin
                        if (timer == 0) begin
                            waddr_packet <= `RST_ADDR;
                            wdata_packet <= 1; 
                            {waddr_valid_packet, wdata_valid_packet} <= 3;
                            timer <= 1;
                        end else begin
                            if (tl.sys.rst) begin
                                timer <= 0;
                                testState <= CHECK;
                            end
                        end
                    end
                    // Read from MAX_ILA address
                    if (test_num == 1) begin
                        if (timer == 0) begin
                            raddr_packet <= `MAX_BURST_SIZE_ADDR;
                            raddr_valid_packet <= 1; 
                            timer <= 1;
                        end else begin
                            if (rdata_valid_out && ps_read_rdy) begin
                                timer <= 0;
                                testState <= CHECK;
                            end
                        end
                    end
                    //Send long pwl wave 
                    if (test_num == 2) begin
                        if (timer < 7) timer <= timer + 1;
                        else begin
                            if (periods == PERIODS_TO_CHECK) begin
                                testState <= CHECK;
                                timer <= 0; 
                            end
                        end

                        if (timer == 0) begin
                            waddr_packet <= `PWL_PREP_ADDR;
                            wdata_packet <= 1; 
                            {waddr_valid_packet, wdata_valid_packet} <= 3;
                            testState <= WRESP; 
                        end 
                        if (timer == 5) send_dma_buff <= 1;                        
                    end
                end
                WRESP: begin
                    if (wresp_valid_out && ps_wresp_rdy) begin
                        if (wresp_out != `OKAY) begin
                            kill_tb <= 1; 
                            testState <= DONE; 
                        end else testState <= TEST; 
                    end
                end 
                CHECK: begin
                    test_num <= test_num + 1;
                    testState <= (test_num < TOTAL_TESTS-1)? TEST : DONE; 
                end 

                DONE: begin 
                    done <= {testsFailed == 0 && ~kill_tb,1'b1}; 
                    testState <= IDLE; 
                    test_num <= 0; 
                end 
            endcase
            if (waddr_valid_packet) waddr_valid_packet <= 0; 
            if (wdata_valid_packet) wdata_valid_packet <= 0; 
            if (raddr_valid_packet) raddr_valid_packet <= 0; 

            if (test_num == 2) begin
                if (test_check[0]) begin
                    if (test_check[1]) begin 
                        testsPassed <= testsPassed + 1;
                        if (VERBOSE) $write("%c[1;32m",27); 
                        if (VERBOSE) $write("t%0d_%0d+ ",test_num,exp_i);
                        if (VERBOSE) $write("%c[0m",27); 
                    end 
                    else begin 
                        testsFailed <= testsFailed + 1; 
                        if (VERBOSE) $write("%c[1;31m",27); 
                        if (VERBOSE) $write("t%0d_%0d- ",test_num,exp_i);
                        if (VERBOSE) $write("%c[0m",27); 
                    end 
                    if (VERBOSE && checked_full_wave) $write("\nChecked period #%0d\n",periods+1);
                end 
            end else begin
                if (test_check[0]) begin
                    if (test_check[1]) begin 
                        testsPassed <= testsPassed + 1;
                        if (VERBOSE) $write("%c[1;32m",27); 
                        if (VERBOSE) $write("t%0d+ ",test_num);
                        if (VERBOSE) $write("%c[0m",27); 
                    end 
                    else begin 
                        testsFailed <= testsFailed + 1; 
                        if (VERBOSE) $write("%c[1;31m",27); 
                        if (VERBOSE) $write("t%0d- ",test_num);
                        if (VERBOSE) $write("%c[0m",27); 
                    end 
                end 
            end

        end
    end

    logic[1:0] testNum_edge, new_sample_edge;
    logic go; 
    enum logic {WATCH, PANIC} panicState; 
    logic[$clog2(TIMEOUT):0] timeout_cntr; 
    edetect testNum_edetect(.clk(clk), .rst(rst),
                            .val(test_num+exp_i),
                            .comb_posedge_out(testNum_edge)); 

    always_ff @(posedge clk) begin 
        if (rst) begin 
            {timeout_cntr,panic} <= 0;
            panicState <= WATCH;
            go <= 0; 
        end 
        else begin
            if (go) begin
                case(panicState) 
                    WATCH: begin
                        if (timeout_cntr <= TIMEOUT) begin
                            if (testNum_edge == 1) timeout_cntr <= 0;
                            else timeout_cntr <= timeout_cntr + 1;
                        end else begin
                            panic <= 1; 
                            panicState <= PANIC; 
                        end 
                    end 
                    PANIC: if (panic) panic <= 0; 
                endcase
            end 
            if (start) go <= 1; 
        end
    end 

    always begin
        #5;  
        clk = !clk;
    end
     
    initial begin
        clk = 0;
        rst = 0; 
        `flash_sig(rst); 
        while (~start) #1; 
        if (VERBOSE) $display("\n############ Starting Top Test ############");
        #100;
        while (testState != DONE && timeout_cntr < TIMEOUT) #10;
        if (timeout_cntr < TIMEOUT) begin
            if (testsFailed != 0) begin 
                if (VERBOSE) $write("%c[1;31m",27); 
                if (VERBOSE) $display("\nTop Tests Failed :((\n");
                if (VERBOSE) $write("%c[0m",27);
            end else begin 
                if (VERBOSE) $write("%c[1;32m",27); 
                if (VERBOSE) $display("\nTop Tests Passed :))\n");
                if (VERBOSE) $write("%c[0m",27); 
            end
            #100;
        end else begin
            $write("%c[1;31m",27); 
            $display("\nTop Tests Timed out on test %d!\n", test_num);
            $write("%c[0m",27);
            #100; 
        end
    end 

endmodule 

`default_nettype wire
