`default_nettype none
`timescale 1ns / 1ps
import mem_layout_pkg::*;

module pwl2_tb();
    localparam SAMPLE_WIDTH = 16;
    localparam BATCH_WIDTH = 48; 
    localparam NSAMPLES = BATCH_WIDTH/SAMPLE_WIDTH; 
    localparam NUM_OF_POINTS = 35; 

    logic clk,rst;
    logic[`MEM_SIZE-1:0] fresh_bits; 
    logic[`BATCH_WIDTH-1:0] dac_batch; 
    logic[`BATCH_SAMPLES-1:0][`SAMPLE_WIDTH-1:0] dac_samples; 
    logic[1:0] valid_dac_edge; 
    logic dac0_rdy, valid_dac_batch; 
    logic[7:0] timer; 
    logic[NUM_OF_POINTS-1:0][`DMA_DATA_WIDTH-1:0] dma_buff;
    logic[`PWL_BRAM_DEPTH-1:0][`BATCH_SAMPLES-1:0][`SAMPLE_WIDTH-1:0] expected_batches;
    logic[`BATCH_SAMPLES-1:0][`SAMPLE_WIDTH-1:0] curr_expected_batch;
    logic[$clog2(`PWL_BRAM_DEPTH):0] exp_i; 
    enum logic[1:0] {IDLE, SEND, CHECK} testState; 
    logic[31:0] correct_vals;
    logic[1:0] correct_edge; 
    Axis_IF #(`DMA_DATA_WIDTH) pwl_dma_if(); 

    assign dac0_rdy = 1; 
    assign curr_expected_batch = expected_batches[exp_i];
    //DMA BUFFER TO SEND
    assign dma_buff = {48'h744000000000, 48'h70de11bffffb, 48'h6c5010350001, 48'h67d40eac0001, 48'h63460d360001, 48'h5ecb0bad0001, 48'h5a3c0a240001, 48'h55c108ae0001, 48'h52720d5effff, 48'h509c14d1fffc, 48'h4dd12ba3fff8, 48'h4c7e35dafff8, 48'h4b3f3ffffff8, 48'h4a7032db0010, 48'h484e2cca0003, 48'h463f26cc0003, 48'h43291b800004, 48'h408414be0003, 48'h3ddf0dfb0003, 48'h3836089a0001, 48'h3755105dfff7, 48'h364d18a9fff8, 48'h35dc201dffef, 48'h35592790fff1, 48'h31162dddffff, 48'h29cf2d400001, 48'h22892ca20001, 48'h1bec2b540001, 48'h1b432c19ffff, 48'h1b3012830159, 48'h1aac00000024, 48'h13fc0076ffff, 48'hd4c00ecffff, 48'h6af014effff, 48'h1};
    //EXPECTED OUTPUT
    assign expected_batches = {0,{16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000},
                                {16'h00da, 16'h00df, 16'h00e4, 16'h00e9, 16'h00ee, 16'h00f3, 16'h00f8, 16'h00fd, 16'h0102, 16'h0107, 16'h010c, 16'h0111, 16'h0116, 16'h011b, 16'h0120, 16'h0125, 16'h012a, 16'h012f, 16'h0134, 16'h0139, 16'h013e, 16'h0143, 16'h0148, 16'h014d, 16'h0152, 16'h0157, 16'h015c, 16'h0161, 16'h0166, 16'h016b, 16'h0170, 16'h0175, 16'h017a, 16'h017f, 16'h0184, 16'h0189, 16'h018e, 16'h0193, 16'h0198, 16'h019d, 16'h01a2, 16'h01a7, 16'h01ac, 16'h01b1, 16'h01b6, 16'h01bb, 16'h01c0, 16'h01c5, 16'h01ca, 16'h01cf, 16'h01d4, 16'h01d9, 16'h01de, 16'h01e3, 16'h01e8, 16'h01ed, 16'h01f2, 16'h01f7, 16'h01fc, 16'h0201, 16'h0206, 16'h020b, 16'h0210, 16'h0215},
                                {16'h021a, 16'h021f, 16'h0224, 16'h0229, 16'h022e, 16'h0233, 16'h0238, 16'h023d, 16'h0242, 16'h0247, 16'h024c, 16'h0251, 16'h0256, 16'h025b, 16'h0260, 16'h0265, 16'h026a, 16'h026f, 16'h0274, 16'h0279, 16'h027e, 16'h0283, 16'h0288, 16'h028d, 16'h0292, 16'h0297, 16'h029c, 16'h02a1, 16'h02a6, 16'h02ab, 16'h02b0, 16'h02b5, 16'h02ba, 16'h02bf, 16'h02c4, 16'h02c9, 16'h02ce, 16'h02d3, 16'h02d8, 16'h02dd, 16'h02e2, 16'h02e7, 16'h02ec, 16'h02f1, 16'h02f6, 16'h02fb, 16'h0300, 16'h0305, 16'h030a, 16'h030f, 16'h0314, 16'h0319, 16'h031e, 16'h0323, 16'h0328, 16'h032d, 16'h0332, 16'h0337, 16'h033c, 16'h0341, 16'h0346, 16'h034b, 16'h0350, 16'h0355},
                                {16'h035a, 16'h035f, 16'h0364, 16'h0369, 16'h036e, 16'h0373, 16'h0378, 16'h037d, 16'h0382, 16'h0387, 16'h038c, 16'h0391, 16'h0396, 16'h039b, 16'h03a0, 16'h03a5, 16'h03aa, 16'h03af, 16'h03b4, 16'h03b9, 16'h03be, 16'h03c3, 16'h03c8, 16'h03cd, 16'h03d2, 16'h03d7, 16'h03dc, 16'h03e1, 16'h03e6, 16'h03eb, 16'h03f0, 16'h03f5, 16'h03fa, 16'h03ff, 16'h0404, 16'h0409, 16'h040e, 16'h0413, 16'h0418, 16'h041d, 16'h0422, 16'h0427, 16'h042c, 16'h0431, 16'h0436, 16'h043b, 16'h0440, 16'h0445, 16'h044a, 16'h044f, 16'h0454, 16'h0459, 16'h045e, 16'h0463, 16'h0468, 16'h046d, 16'h0472, 16'h0477, 16'h047c, 16'h0481, 16'h0486, 16'h048b, 16'h0490, 16'h0495},
                                {16'h049a, 16'h049f, 16'h04a4, 16'h04a9, 16'h04ae, 16'h04b3, 16'h04b8, 16'h04bd, 16'h04c2, 16'h04c7, 16'h04cc, 16'h04d1, 16'h04d6, 16'h04db, 16'h04e0, 16'h04e5, 16'h04ea, 16'h04ef, 16'h04f4, 16'h04f9, 16'h04fe, 16'h0503, 16'h0508, 16'h050d, 16'h0512, 16'h0517, 16'h051c, 16'h0521, 16'h0526, 16'h052b, 16'h0530, 16'h0535, 16'h053a, 16'h053f, 16'h0544, 16'h0549, 16'h054e, 16'h0553, 16'h0558, 16'h055d, 16'h0562, 16'h0567, 16'h056c, 16'h0571, 16'h0576, 16'h057b, 16'h0580, 16'h0585, 16'h058a, 16'h058f, 16'h0594, 16'h0599, 16'h059e, 16'h05a3, 16'h05a8, 16'h05ad, 16'h05b2, 16'h05b7, 16'h05bc, 16'h05c1, 16'h05c6, 16'h05cb, 16'h05d0, 16'h05d5},
                                {16'h05da, 16'h05df, 16'h05e4, 16'h05e9, 16'h05ee, 16'h05f3, 16'h05f8, 16'h05fd, 16'h0602, 16'h0607, 16'h060c, 16'h0611, 16'h0616, 16'h061b, 16'h0620, 16'h0625, 16'h062a, 16'h062f, 16'h0634, 16'h0639, 16'h063e, 16'h0643, 16'h0648, 16'h064d, 16'h0652, 16'h0657, 16'h065c, 16'h0661, 16'h0666, 16'h066b, 16'h0670, 16'h0675, 16'h067a, 16'h067f, 16'h0684, 16'h0689, 16'h068e, 16'h0693, 16'h0698, 16'h069d, 16'h06a2, 16'h06a7, 16'h06ac, 16'h06b1, 16'h06b6, 16'h06bb, 16'h06c0, 16'h06c5, 16'h06ca, 16'h06cf, 16'h06d4, 16'h06d9, 16'h06de, 16'h06e3, 16'h06e8, 16'h06ed, 16'h06f2, 16'h06f7, 16'h06fc, 16'h0701, 16'h0706, 16'h070b, 16'h0710, 16'h0715},
                                {16'h071a, 16'h071f, 16'h0724, 16'h0729, 16'h072e, 16'h0733, 16'h0738, 16'h073d, 16'h0742, 16'h0747, 16'h074c, 16'h0751, 16'h0756, 16'h075b, 16'h0760, 16'h0765, 16'h076a, 16'h076f, 16'h0774, 16'h0779, 16'h077e, 16'h0783, 16'h0788, 16'h078d, 16'h0792, 16'h0797, 16'h079c, 16'h07a1, 16'h07a6, 16'h07ab, 16'h07b0, 16'h07b5, 16'h07ba, 16'h07bf, 16'h07c4, 16'h07c9, 16'h07ce, 16'h07d3, 16'h07d8, 16'h07dd, 16'h07e2, 16'h07e7, 16'h07ec, 16'h07f1, 16'h07f6, 16'h07fb, 16'h0800, 16'h0805, 16'h080a, 16'h080f, 16'h0814, 16'h0819, 16'h081e, 16'h0823, 16'h0828, 16'h082d, 16'h0832, 16'h0837, 16'h083c, 16'h0841, 16'h0846, 16'h084b, 16'h0850, 16'h0855},
                                {16'h085a, 16'h085f, 16'h0864, 16'h0869, 16'h086e, 16'h0873, 16'h0878, 16'h087d, 16'h0882, 16'h0887, 16'h088c, 16'h0891, 16'h0896, 16'h089b, 16'h08a0, 16'h08a5, 16'h08aa, 16'h08af, 16'h08b4, 16'h08b9, 16'h08be, 16'h08c3, 16'h08c8, 16'h08cd, 16'h08d2, 16'h08d7, 16'h08dc, 16'h08e1, 16'h08e6, 16'h08eb, 16'h08f0, 16'h08f5, 16'h08fa, 16'h08ff, 16'h0904, 16'h0909, 16'h090e, 16'h0913, 16'h0918, 16'h091d, 16'h0922, 16'h0927, 16'h092c, 16'h0931, 16'h0936, 16'h093b, 16'h0940, 16'h0945, 16'h094a, 16'h094f, 16'h0954, 16'h0959, 16'h095e, 16'h0963, 16'h0968, 16'h096d, 16'h0972, 16'h0977, 16'h097c, 16'h0981, 16'h0986, 16'h098b, 16'h0990, 16'h0995},
                                {16'h099a, 16'h099f, 16'h09a4, 16'h09a9, 16'h09ae, 16'h09b3, 16'h09b8, 16'h09bd, 16'h09c2, 16'h09c7, 16'h09cc, 16'h09d1, 16'h09d6, 16'h09db, 16'h09e0, 16'h09e5, 16'h09ea, 16'h09ef, 16'h09f4, 16'h09f9, 16'h09fe, 16'h0a03, 16'h0a08, 16'h0a0d, 16'h0a12, 16'h0a17, 16'h0a1c, 16'h0a21, 16'h0a26, 16'h0a2b, 16'h0a30, 16'h0a35, 16'h0a3a, 16'h0a3f, 16'h0a44, 16'h0a49, 16'h0a4e, 16'h0a53, 16'h0a58, 16'h0a5d, 16'h0a62, 16'h0a67, 16'h0a6c, 16'h0a71, 16'h0a76, 16'h0a7b, 16'h0a80, 16'h0a85, 16'h0a8a, 16'h0a8f, 16'h0a94, 16'h0a99, 16'h0a9e, 16'h0aa3, 16'h0aa8, 16'h0aad, 16'h0ab2, 16'h0ab7, 16'h0abc, 16'h0ac1, 16'h0ac6, 16'h0acb, 16'h0ad0, 16'h0ad5},
                                {16'h0ada, 16'h0adf, 16'h0ae4, 16'h0ae9, 16'h0aee, 16'h0af3, 16'h0af8, 16'h0afd, 16'h0b02, 16'h0b07, 16'h0b0c, 16'h0b11, 16'h0b16, 16'h0b1b, 16'h0b20, 16'h0b25, 16'h0b2a, 16'h0b2f, 16'h0b34, 16'h0b39, 16'h0b3e, 16'h0b43, 16'h0b48, 16'h0b4d, 16'h0b52, 16'h0b57, 16'h0b5c, 16'h0b61, 16'h0b66, 16'h0b6b, 16'h0b70, 16'h0b75, 16'h0b7a, 16'h0b7f, 16'h0b84, 16'h0b89, 16'h0b8e, 16'h0b93, 16'h0b98, 16'h0b9d, 16'h0ba2, 16'h0ba7, 16'h0bac, 16'h0bb1, 16'h0bb6, 16'h0bbb, 16'h0bc0, 16'h0bc5, 16'h0bca, 16'h0bcf, 16'h0bd4, 16'h0bd9, 16'h0bde, 16'h0be3, 16'h0be8, 16'h0bed, 16'h0bf2, 16'h0bf7, 16'h0bfc, 16'h0c01, 16'h0c06, 16'h0c0b, 16'h0c10, 16'h0c15},
                                {16'h0c1a, 16'h0c1f, 16'h0c24, 16'h0c29, 16'h0c2e, 16'h0c33, 16'h0c38, 16'h0c3d, 16'h0c42, 16'h0c47, 16'h0c4c, 16'h0c51, 16'h0c56, 16'h0c5b, 16'h0c60, 16'h0c65, 16'h0c6a, 16'h0c6f, 16'h0c74, 16'h0c79, 16'h0c7e, 16'h0c83, 16'h0c88, 16'h0c8d, 16'h0c92, 16'h0c97, 16'h0c9c, 16'h0ca1, 16'h0ca6, 16'h0cab, 16'h0cb0, 16'h0cb5, 16'h0cba, 16'h0cbf, 16'h0cc4, 16'h0cc9, 16'h0cce, 16'h0cd3, 16'h0cd8, 16'h0cdd, 16'h0ce2, 16'h0ce7, 16'h0cec, 16'h0cf1, 16'h0cf6, 16'h0cfb, 16'h0d00, 16'h0d05, 16'h0d0a, 16'h0d0f, 16'h0d14, 16'h0d19, 16'h0d1e, 16'h0d23, 16'h0d28, 16'h0d2d, 16'h0d32, 16'h0d37, 16'h0d3c, 16'h0d41, 16'h0d46, 16'h0d4b, 16'h0d50, 16'h0d55},
                                {16'h0d5a, 16'h0d5f, 16'h0d64, 16'h0d69, 16'h0d6e, 16'h0d73, 16'h0d78, 16'h0d7d, 16'h0d82, 16'h0d87, 16'h0d8c, 16'h0d91, 16'h0d96, 16'h0d9b, 16'h0da0, 16'h0da5, 16'h0daa, 16'h0daf, 16'h0db4, 16'h0db9, 16'h0dbe, 16'h0dc3, 16'h0dc8, 16'h0dcd, 16'h0dd2, 16'h0dd7, 16'h0ddc, 16'h0de1, 16'h0de6, 16'h0deb, 16'h0df0, 16'h0df5, 16'h0dfa, 16'h0dff, 16'h0e04, 16'h0e09, 16'h0e0e, 16'h0e13, 16'h0e18, 16'h0e1d, 16'h0e22, 16'h0e27, 16'h0e2c, 16'h0e31, 16'h0e36, 16'h0e3b, 16'h0e40, 16'h0e45, 16'h0e4a, 16'h0e4f, 16'h0e54, 16'h0e59, 16'h0e5e, 16'h0e63, 16'h0e68, 16'h0e6d, 16'h0e72, 16'h0e77, 16'h0e7c, 16'h0e81, 16'h0e86, 16'h0e8b, 16'h0e90, 16'h0e95},
                                {16'h0e9a, 16'h0e9f, 16'h0ea4, 16'h0ea9, 16'h0eae, 16'h0eb3, 16'h0eb8, 16'h0ebd, 16'h0ec2, 16'h0ec7, 16'h0ecc, 16'h0ed1, 16'h0ed6, 16'h0edb, 16'h0ee0, 16'h0ee5, 16'h0eea, 16'h0eef, 16'h0ef4, 16'h0ef9, 16'h0efe, 16'h0f03, 16'h0f08, 16'h0f0d, 16'h0f12, 16'h0f17, 16'h0f1c, 16'h0f21, 16'h0f26, 16'h0f2b, 16'h0f30, 16'h0f35, 16'h0f3a, 16'h0f3f, 16'h0f44, 16'h0f49, 16'h0f4e, 16'h0f53, 16'h0f58, 16'h0f5d, 16'h0f62, 16'h0f67, 16'h0f6c, 16'h0f71, 16'h0f76, 16'h0f7b, 16'h0f80, 16'h0f85, 16'h0f8a, 16'h0f8f, 16'h0f94, 16'h0f99, 16'h0f9e, 16'h0fa3, 16'h0fa8, 16'h0fad, 16'h0fb2, 16'h0fb7, 16'h0fbc, 16'h0fc1, 16'h0fc6, 16'h0fcb, 16'h0fd0, 16'h0fd5},
                                {16'h0fda, 16'h0fdf, 16'h0fe4, 16'h0fe9, 16'h0fee, 16'h0ff3, 16'h0ff8, 16'h0ffd, 16'h1002, 16'h1007, 16'h100c, 16'h1011, 16'h1016, 16'h101b, 16'h1020, 16'h1025, 16'h102a, 16'h102f, 16'h1034, 16'h1039, 16'h103e, 16'h1043, 16'h1048, 16'h104d, 16'h1052, 16'h1057, 16'h105c, 16'h1061, 16'h1066, 16'h106b, 16'h1070, 16'h1075, 16'h107a, 16'h107f, 16'h1084, 16'h1089, 16'h108e, 16'h1093, 16'h1098, 16'h109d, 16'h10a2, 16'h10a7, 16'h10ac, 16'h10b1, 16'h10b6, 16'h10bb, 16'h10c0, 16'h10c5, 16'h10ca, 16'h10cf, 16'h10d4, 16'h10d9, 16'h10de, 16'h10e3, 16'h10e8, 16'h10ed, 16'h10f2, 16'h10f7, 16'h10fc, 16'h1101, 16'h1106, 16'h110b, 16'h1110, 16'h1115},
                                {16'h111a, 16'h111f, 16'h1124, 16'h1129, 16'h112e, 16'h1133, 16'h1138, 16'h113d, 16'h1142, 16'h1147, 16'h114c, 16'h1151, 16'h1156, 16'h115b, 16'h1160, 16'h1165, 16'h116a, 16'h116f, 16'h1174, 16'h1179, 16'h117e, 16'h1183, 16'h1188, 16'h118d, 16'h1192, 16'h1197, 16'h119c, 16'h11a1, 16'h11a6, 16'h11ab, 16'h11b0, 16'h11b5, 16'h11ba, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf},
                                {16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf},
                                {16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf},
                                {16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf},
                                {16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf},
                                {16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf},
                                {16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf},
                                {16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf},
                                {16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf},
                                {16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf},
                                {16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf},
                                {16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf},
                                {16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11bf, 16'h11be, 16'h11bd, 16'h11bc, 16'h11bb, 16'h11ba, 16'h11b9, 16'h11b8, 16'h11b7, 16'h11b6, 16'h11b5, 16'h11b4, 16'h11b3, 16'h11b2, 16'h11b1, 16'h11b0, 16'h11af, 16'h11ae, 16'h11ad, 16'h11ac, 16'h11ab, 16'h11aa, 16'h11a9, 16'h11a8, 16'h11a7, 16'h11a6, 16'h11a5},
                                {16'h11a4, 16'h11a3, 16'h11a2, 16'h11a1, 16'h11a0, 16'h119f, 16'h119e, 16'h119d, 16'h119c, 16'h119b, 16'h119a, 16'h1199, 16'h1198, 16'h1197, 16'h1196, 16'h1195, 16'h1194, 16'h1193, 16'h1192, 16'h1191, 16'h1190, 16'h118f, 16'h118e, 16'h118d, 16'h118c, 16'h118b, 16'h118a, 16'h1189, 16'h1188, 16'h1187, 16'h1186, 16'h1185, 16'h1184, 16'h1183, 16'h1182, 16'h1181, 16'h1180, 16'h117f, 16'h117e, 16'h117d, 16'h117c, 16'h117b, 16'h117a, 16'h1179, 16'h1178, 16'h1177, 16'h1176, 16'h1175, 16'h1174, 16'h1173, 16'h1172, 16'h1171, 16'h1170, 16'h116f, 16'h116e, 16'h116d, 16'h116c, 16'h116b, 16'h116a, 16'h1169, 16'h1168, 16'h1167, 16'h1166, 16'h1165},
                                {16'h1164, 16'h1163, 16'h1162, 16'h1161, 16'h1160, 16'h115f, 16'h115e, 16'h115d, 16'h115c, 16'h115b, 16'h115a, 16'h1159, 16'h1158, 16'h1157, 16'h1156, 16'h1155, 16'h1154, 16'h1153, 16'h1152, 16'h1151, 16'h1150, 16'h114f, 16'h114e, 16'h114d, 16'h114c, 16'h114b, 16'h114a, 16'h1149, 16'h1148, 16'h1147, 16'h1146, 16'h1145, 16'h1144, 16'h1143, 16'h1142, 16'h1141, 16'h1140, 16'h113f, 16'h113e, 16'h113d, 16'h113c, 16'h113b, 16'h113a, 16'h1139, 16'h1138, 16'h1137, 16'h1136, 16'h1135, 16'h1134, 16'h1133, 16'h1132, 16'h1131, 16'h1130, 16'h112f, 16'h112e, 16'h112d, 16'h112c, 16'h112b, 16'h112a, 16'h1129, 16'h1128, 16'h1127, 16'h1126, 16'h1125},
                                {16'h1124, 16'h1123, 16'h1122, 16'h1121, 16'h1120, 16'h111f, 16'h111e, 16'h111d, 16'h111c, 16'h111b, 16'h111a, 16'h1119, 16'h1118, 16'h1117, 16'h1116, 16'h1115, 16'h1114, 16'h1113, 16'h1112, 16'h1111, 16'h1110, 16'h110f, 16'h110e, 16'h110d, 16'h110c, 16'h110b, 16'h110a, 16'h1109, 16'h1108, 16'h1107, 16'h1106, 16'h1105, 16'h1104, 16'h1103, 16'h1102, 16'h1101, 16'h1100, 16'h10ff, 16'h10fe, 16'h10fd, 16'h10fc, 16'h10fb, 16'h10fa, 16'h10f9, 16'h10f8, 16'h10f7, 16'h10f6, 16'h10f5, 16'h10f4, 16'h10f3, 16'h10f2, 16'h10f1, 16'h10f0, 16'h10ef, 16'h10ee, 16'h10ed, 16'h10ec, 16'h10eb, 16'h10ea, 16'h10e9, 16'h10e8, 16'h10e7, 16'h10e6, 16'h10e5},
                                {16'h10e4, 16'h10e3, 16'h10e2, 16'h10e1, 16'h10e0, 16'h10df, 16'h10de, 16'h10dd, 16'h10dc, 16'h10db, 16'h10da, 16'h10d9, 16'h10d8, 16'h10d7, 16'h10d6, 16'h10d5, 16'h10d4, 16'h10d3, 16'h10d2, 16'h10d1, 16'h10d0, 16'h10cf, 16'h10ce, 16'h10cd, 16'h10cc, 16'h10cb, 16'h10ca, 16'h10c9, 16'h10c8, 16'h10c7, 16'h10c6, 16'h10c5, 16'h10c4, 16'h10c3, 16'h10c2, 16'h10c1, 16'h10c0, 16'h10bf, 16'h10be, 16'h10bd, 16'h10bc, 16'h10bb, 16'h10ba, 16'h10b9, 16'h10b8, 16'h10b7, 16'h10b6, 16'h10b5, 16'h10b4, 16'h10b3, 16'h10b2, 16'h10b1, 16'h10b0, 16'h10af, 16'h10ae, 16'h10ad, 16'h10ac, 16'h10ab, 16'h10aa, 16'h10a9, 16'h10a8, 16'h10a7, 16'h10a6, 16'h10a5},
                                {16'h10a4, 16'h10a3, 16'h10a2, 16'h10a1, 16'h10a0, 16'h109f, 16'h109e, 16'h109d, 16'h109c, 16'h109b, 16'h109a, 16'h1099, 16'h1098, 16'h1097, 16'h1096, 16'h1095, 16'h1094, 16'h1093, 16'h1092, 16'h1091, 16'h1090, 16'h108f, 16'h108e, 16'h108d, 16'h108c, 16'h108b, 16'h108a, 16'h1089, 16'h1088, 16'h1087, 16'h1086, 16'h1085, 16'h1084, 16'h1083, 16'h1082, 16'h1081, 16'h1080, 16'h107f, 16'h107e, 16'h107d, 16'h107c, 16'h107b, 16'h107a, 16'h1079, 16'h1078, 16'h1077, 16'h1076, 16'h1075, 16'h1074, 16'h1073, 16'h1072, 16'h1071, 16'h1070, 16'h106f, 16'h106e, 16'h106d, 16'h106c, 16'h106b, 16'h106a, 16'h1069, 16'h1068, 16'h1067, 16'h1066, 16'h1065},
                                {16'h1064, 16'h1063, 16'h1062, 16'h1061, 16'h1060, 16'h105f, 16'h105e, 16'h105d, 16'h105c, 16'h105b, 16'h105a, 16'h1059, 16'h1058, 16'h1057, 16'h1056, 16'h1055, 16'h1054, 16'h1053, 16'h1052, 16'h1051, 16'h1050, 16'h104f, 16'h104e, 16'h104d, 16'h104c, 16'h104b, 16'h104a, 16'h1049, 16'h1048, 16'h1047, 16'h1046, 16'h1045, 16'h1044, 16'h1043, 16'h1042, 16'h1041, 16'h1040, 16'h103f, 16'h103e, 16'h103d, 16'h103c, 16'h103b, 16'h103a, 16'h1039, 16'h1038, 16'h1037, 16'h1036, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035},
                                {16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035},
                                {16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035},
                                {16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035},
                                {16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035},
                                {16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035},
                                {16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035},
                                {16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035},
                                {16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035},
                                {16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035},
                                {16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035},
                                {16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035},
                                {16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1035, 16'h1034, 16'h1033, 16'h1032, 16'h1031, 16'h1030, 16'h102f, 16'h102e, 16'h102d, 16'h102c, 16'h102b, 16'h102a, 16'h1029, 16'h1028, 16'h1027, 16'h1026, 16'h1025, 16'h1024, 16'h1023, 16'h1022, 16'h1021, 16'h1020, 16'h101f, 16'h101e, 16'h101d, 16'h101c, 16'h101b, 16'h101a, 16'h1019, 16'h1018},
                                {16'h1017, 16'h1016, 16'h1015, 16'h1014, 16'h1013, 16'h1012, 16'h1011, 16'h1010, 16'h100f, 16'h100e, 16'h100d, 16'h100c, 16'h100b, 16'h100a, 16'h1009, 16'h1008, 16'h1007, 16'h1006, 16'h1005, 16'h1004, 16'h1003, 16'h1002, 16'h1001, 16'h1000, 16'h0fff, 16'h0ffe, 16'h0ffd, 16'h0ffc, 16'h0ffb, 16'h0ffa, 16'h0ff9, 16'h0ff8, 16'h0ff7, 16'h0ff6, 16'h0ff5, 16'h0ff4, 16'h0ff3, 16'h0ff2, 16'h0ff1, 16'h0ff0, 16'h0fef, 16'h0fee, 16'h0fed, 16'h0fec, 16'h0feb, 16'h0fea, 16'h0fe9, 16'h0fe8, 16'h0fe7, 16'h0fe6, 16'h0fe5, 16'h0fe4, 16'h0fe3, 16'h0fe2, 16'h0fe1, 16'h0fe0, 16'h0fdf, 16'h0fde, 16'h0fdd, 16'h0fdc, 16'h0fdb, 16'h0fda, 16'h0fd9, 16'h0fd8},
                                {16'h0fd7, 16'h0fd6, 16'h0fd5, 16'h0fd4, 16'h0fd3, 16'h0fd2, 16'h0fd1, 16'h0fd0, 16'h0fcf, 16'h0fce, 16'h0fcd, 16'h0fcc, 16'h0fcb, 16'h0fca, 16'h0fc9, 16'h0fc8, 16'h0fc7, 16'h0fc6, 16'h0fc5, 16'h0fc4, 16'h0fc3, 16'h0fc2, 16'h0fc1, 16'h0fc0, 16'h0fbf, 16'h0fbe, 16'h0fbd, 16'h0fbc, 16'h0fbb, 16'h0fba, 16'h0fb9, 16'h0fb8, 16'h0fb7, 16'h0fb6, 16'h0fb5, 16'h0fb4, 16'h0fb3, 16'h0fb2, 16'h0fb1, 16'h0fb0, 16'h0faf, 16'h0fae, 16'h0fad, 16'h0fac, 16'h0fab, 16'h0faa, 16'h0fa9, 16'h0fa8, 16'h0fa7, 16'h0fa6, 16'h0fa5, 16'h0fa4, 16'h0fa3, 16'h0fa2, 16'h0fa1, 16'h0fa0, 16'h0f9f, 16'h0f9e, 16'h0f9d, 16'h0f9c, 16'h0f9b, 16'h0f9a, 16'h0f99, 16'h0f98},
                                {16'h0f97, 16'h0f96, 16'h0f95, 16'h0f94, 16'h0f93, 16'h0f92, 16'h0f91, 16'h0f90, 16'h0f8f, 16'h0f8e, 16'h0f8d, 16'h0f8c, 16'h0f8b, 16'h0f8a, 16'h0f89, 16'h0f88, 16'h0f87, 16'h0f86, 16'h0f85, 16'h0f84, 16'h0f83, 16'h0f82, 16'h0f81, 16'h0f80, 16'h0f7f, 16'h0f7e, 16'h0f7d, 16'h0f7c, 16'h0f7b, 16'h0f7a, 16'h0f79, 16'h0f78, 16'h0f77, 16'h0f76, 16'h0f75, 16'h0f74, 16'h0f73, 16'h0f72, 16'h0f71, 16'h0f70, 16'h0f6f, 16'h0f6e, 16'h0f6d, 16'h0f6c, 16'h0f6b, 16'h0f6a, 16'h0f69, 16'h0f68, 16'h0f67, 16'h0f66, 16'h0f65, 16'h0f64, 16'h0f63, 16'h0f62, 16'h0f61, 16'h0f60, 16'h0f5f, 16'h0f5e, 16'h0f5d, 16'h0f5c, 16'h0f5b, 16'h0f5a, 16'h0f59, 16'h0f58},
                                {16'h0f57, 16'h0f56, 16'h0f55, 16'h0f54, 16'h0f53, 16'h0f52, 16'h0f51, 16'h0f50, 16'h0f4f, 16'h0f4e, 16'h0f4d, 16'h0f4c, 16'h0f4b, 16'h0f4a, 16'h0f49, 16'h0f48, 16'h0f47, 16'h0f46, 16'h0f45, 16'h0f44, 16'h0f43, 16'h0f42, 16'h0f41, 16'h0f40, 16'h0f3f, 16'h0f3e, 16'h0f3d, 16'h0f3c, 16'h0f3b, 16'h0f3a, 16'h0f39, 16'h0f38, 16'h0f37, 16'h0f36, 16'h0f35, 16'h0f34, 16'h0f33, 16'h0f32, 16'h0f31, 16'h0f30, 16'h0f2f, 16'h0f2e, 16'h0f2d, 16'h0f2c, 16'h0f2b, 16'h0f2a, 16'h0f29, 16'h0f28, 16'h0f27, 16'h0f26, 16'h0f25, 16'h0f24, 16'h0f23, 16'h0f22, 16'h0f21, 16'h0f20, 16'h0f1f, 16'h0f1e, 16'h0f1d, 16'h0f1c, 16'h0f1b, 16'h0f1a, 16'h0f19, 16'h0f18},
                                {16'h0f17, 16'h0f16, 16'h0f15, 16'h0f14, 16'h0f13, 16'h0f12, 16'h0f11, 16'h0f10, 16'h0f0f, 16'h0f0e, 16'h0f0d, 16'h0f0c, 16'h0f0b, 16'h0f0a, 16'h0f09, 16'h0f08, 16'h0f07, 16'h0f06, 16'h0f05, 16'h0f04, 16'h0f03, 16'h0f02, 16'h0f01, 16'h0f00, 16'h0eff, 16'h0efe, 16'h0efd, 16'h0efc, 16'h0efb, 16'h0efa, 16'h0ef9, 16'h0ef8, 16'h0ef7, 16'h0ef6, 16'h0ef5, 16'h0ef4, 16'h0ef3, 16'h0ef2, 16'h0ef1, 16'h0ef0, 16'h0eef, 16'h0eee, 16'h0eed, 16'h0eec, 16'h0eeb, 16'h0eea, 16'h0ee9, 16'h0ee8, 16'h0ee7, 16'h0ee6, 16'h0ee5, 16'h0ee4, 16'h0ee3, 16'h0ee2, 16'h0ee1, 16'h0ee0, 16'h0edf, 16'h0ede, 16'h0edd, 16'h0edc, 16'h0edb, 16'h0eda, 16'h0ed9, 16'h0ed8},
                                {16'h0ed7, 16'h0ed6, 16'h0ed5, 16'h0ed4, 16'h0ed3, 16'h0ed2, 16'h0ed1, 16'h0ed0, 16'h0ecf, 16'h0ece, 16'h0ecd, 16'h0ecc, 16'h0ecb, 16'h0eca, 16'h0ec9, 16'h0ec8, 16'h0ec7, 16'h0ec6, 16'h0ec5, 16'h0ec4, 16'h0ec3, 16'h0ec2, 16'h0ec1, 16'h0ec0, 16'h0ebf, 16'h0ebe, 16'h0ebd, 16'h0ebc, 16'h0ebb, 16'h0eba, 16'h0eb9, 16'h0eb8, 16'h0eb7, 16'h0eb6, 16'h0eb5, 16'h0eb4, 16'h0eb3, 16'h0eb2, 16'h0eb1, 16'h0eb0, 16'h0eaf, 16'h0eae, 16'h0ead, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac},
                                {16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac},
                                {16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac},
                                {16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac},
                                {16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac},
                                {16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac},
                                {16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac},
                                {16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac},
                                {16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac},
                                {16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac},
                                {16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac},
                                {16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac},
                                {16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac},
                                {16'h0eac, 16'h0eac, 16'h0eac, 16'h0eac, 16'h0eab, 16'h0eaa, 16'h0ea9, 16'h0ea8, 16'h0ea7, 16'h0ea6, 16'h0ea5, 16'h0ea4, 16'h0ea3, 16'h0ea2, 16'h0ea1, 16'h0ea0, 16'h0e9f, 16'h0e9e, 16'h0e9d, 16'h0e9c, 16'h0e9b, 16'h0e9a, 16'h0e99, 16'h0e98, 16'h0e97, 16'h0e96, 16'h0e95, 16'h0e94, 16'h0e93, 16'h0e92, 16'h0e91, 16'h0e90, 16'h0e8f, 16'h0e8e, 16'h0e8d, 16'h0e8c, 16'h0e8b, 16'h0e8a, 16'h0e89, 16'h0e88, 16'h0e87, 16'h0e86, 16'h0e85, 16'h0e84, 16'h0e83, 16'h0e82, 16'h0e81, 16'h0e80, 16'h0e7f, 16'h0e7e, 16'h0e7d, 16'h0e7c, 16'h0e7b, 16'h0e7a, 16'h0e79, 16'h0e78, 16'h0e77, 16'h0e76, 16'h0e75, 16'h0e74, 16'h0e73, 16'h0e72, 16'h0e71, 16'h0e70},
                                {16'h0e6f, 16'h0e6e, 16'h0e6d, 16'h0e6c, 16'h0e6b, 16'h0e6a, 16'h0e69, 16'h0e68, 16'h0e67, 16'h0e66, 16'h0e65, 16'h0e64, 16'h0e63, 16'h0e62, 16'h0e61, 16'h0e60, 16'h0e5f, 16'h0e5e, 16'h0e5d, 16'h0e5c, 16'h0e5b, 16'h0e5a, 16'h0e59, 16'h0e58, 16'h0e57, 16'h0e56, 16'h0e55, 16'h0e54, 16'h0e53, 16'h0e52, 16'h0e51, 16'h0e50, 16'h0e4f, 16'h0e4e, 16'h0e4d, 16'h0e4c, 16'h0e4b, 16'h0e4a, 16'h0e49, 16'h0e48, 16'h0e47, 16'h0e46, 16'h0e45, 16'h0e44, 16'h0e43, 16'h0e42, 16'h0e41, 16'h0e40, 16'h0e3f, 16'h0e3e, 16'h0e3d, 16'h0e3c, 16'h0e3b, 16'h0e3a, 16'h0e39, 16'h0e38, 16'h0e37, 16'h0e36, 16'h0e35, 16'h0e34, 16'h0e33, 16'h0e32, 16'h0e31, 16'h0e30},
                                {16'h0e2f, 16'h0e2e, 16'h0e2d, 16'h0e2c, 16'h0e2b, 16'h0e2a, 16'h0e29, 16'h0e28, 16'h0e27, 16'h0e26, 16'h0e25, 16'h0e24, 16'h0e23, 16'h0e22, 16'h0e21, 16'h0e20, 16'h0e1f, 16'h0e1e, 16'h0e1d, 16'h0e1c, 16'h0e1b, 16'h0e1a, 16'h0e19, 16'h0e18, 16'h0e17, 16'h0e16, 16'h0e15, 16'h0e14, 16'h0e13, 16'h0e12, 16'h0e11, 16'h0e10, 16'h0e0f, 16'h0e0e, 16'h0e0d, 16'h0e0c, 16'h0e0b, 16'h0e0a, 16'h0e09, 16'h0e08, 16'h0e07, 16'h0e06, 16'h0e05, 16'h0e04, 16'h0e03, 16'h0e02, 16'h0e01, 16'h0e00, 16'h0dff, 16'h0dfe, 16'h0dfd, 16'h0dfc, 16'h0dfb, 16'h0dfa, 16'h0df9, 16'h0df8, 16'h0df7, 16'h0df6, 16'h0df5, 16'h0df4, 16'h0df3, 16'h0df2, 16'h0df1, 16'h0df0},
                                {16'h0def, 16'h0dee, 16'h0ded, 16'h0dec, 16'h0deb, 16'h0dea, 16'h0de9, 16'h0de8, 16'h0de7, 16'h0de6, 16'h0de5, 16'h0de4, 16'h0de3, 16'h0de2, 16'h0de1, 16'h0de0, 16'h0ddf, 16'h0dde, 16'h0ddd, 16'h0ddc, 16'h0ddb, 16'h0dda, 16'h0dd9, 16'h0dd8, 16'h0dd7, 16'h0dd6, 16'h0dd5, 16'h0dd4, 16'h0dd3, 16'h0dd2, 16'h0dd1, 16'h0dd0, 16'h0dcf, 16'h0dce, 16'h0dcd, 16'h0dcc, 16'h0dcb, 16'h0dca, 16'h0dc9, 16'h0dc8, 16'h0dc7, 16'h0dc6, 16'h0dc5, 16'h0dc4, 16'h0dc3, 16'h0dc2, 16'h0dc1, 16'h0dc0, 16'h0dbf, 16'h0dbe, 16'h0dbd, 16'h0dbc, 16'h0dbb, 16'h0dba, 16'h0db9, 16'h0db8, 16'h0db7, 16'h0db6, 16'h0db5, 16'h0db4, 16'h0db3, 16'h0db2, 16'h0db1, 16'h0db0},
                                {16'h0daf, 16'h0dae, 16'h0dad, 16'h0dac, 16'h0dab, 16'h0daa, 16'h0da9, 16'h0da8, 16'h0da7, 16'h0da6, 16'h0da5, 16'h0da4, 16'h0da3, 16'h0da2, 16'h0da1, 16'h0da0, 16'h0d9f, 16'h0d9e, 16'h0d9d, 16'h0d9c, 16'h0d9b, 16'h0d9a, 16'h0d99, 16'h0d98, 16'h0d97, 16'h0d96, 16'h0d95, 16'h0d94, 16'h0d93, 16'h0d92, 16'h0d91, 16'h0d90, 16'h0d8f, 16'h0d8e, 16'h0d8d, 16'h0d8c, 16'h0d8b, 16'h0d8a, 16'h0d89, 16'h0d88, 16'h0d87, 16'h0d86, 16'h0d85, 16'h0d84, 16'h0d83, 16'h0d82, 16'h0d81, 16'h0d80, 16'h0d7f, 16'h0d7e, 16'h0d7d, 16'h0d7c, 16'h0d7b, 16'h0d7a, 16'h0d79, 16'h0d78, 16'h0d77, 16'h0d76, 16'h0d75, 16'h0d74, 16'h0d73, 16'h0d72, 16'h0d71, 16'h0d70},
                                {16'h0d6f, 16'h0d6e, 16'h0d6d, 16'h0d6c, 16'h0d6b, 16'h0d6a, 16'h0d69, 16'h0d68, 16'h0d67, 16'h0d66, 16'h0d65, 16'h0d64, 16'h0d63, 16'h0d62, 16'h0d61, 16'h0d60, 16'h0d5f, 16'h0d5e, 16'h0d5d, 16'h0d5c, 16'h0d5b, 16'h0d5a, 16'h0d59, 16'h0d58, 16'h0d57, 16'h0d56, 16'h0d55, 16'h0d54, 16'h0d53, 16'h0d52, 16'h0d51, 16'h0d50, 16'h0d4f, 16'h0d4e, 16'h0d4d, 16'h0d4c, 16'h0d4b, 16'h0d4a, 16'h0d49, 16'h0d48, 16'h0d47, 16'h0d46, 16'h0d45, 16'h0d44, 16'h0d43, 16'h0d42, 16'h0d41, 16'h0d40, 16'h0d3f, 16'h0d3e, 16'h0d3d, 16'h0d3c, 16'h0d3b, 16'h0d3a, 16'h0d39, 16'h0d38, 16'h0d37, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36},
                                {16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36},
                                {16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36},
                                {16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36},
                                {16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36},
                                {16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36},
                                {16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36},
                                {16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36},
                                {16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36},
                                {16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36},
                                {16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36},
                                {16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36},
                                {16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d36, 16'h0d35, 16'h0d34, 16'h0d33, 16'h0d32, 16'h0d31, 16'h0d30, 16'h0d2f, 16'h0d2e, 16'h0d2d, 16'h0d2c, 16'h0d2b, 16'h0d2a, 16'h0d29, 16'h0d28, 16'h0d27, 16'h0d26, 16'h0d25, 16'h0d24, 16'h0d23, 16'h0d22},
                                {16'h0d21, 16'h0d20, 16'h0d1f, 16'h0d1e, 16'h0d1d, 16'h0d1c, 16'h0d1b, 16'h0d1a, 16'h0d19, 16'h0d18, 16'h0d17, 16'h0d16, 16'h0d15, 16'h0d14, 16'h0d13, 16'h0d12, 16'h0d11, 16'h0d10, 16'h0d0f, 16'h0d0e, 16'h0d0d, 16'h0d0c, 16'h0d0b, 16'h0d0a, 16'h0d09, 16'h0d08, 16'h0d07, 16'h0d06, 16'h0d05, 16'h0d04, 16'h0d03, 16'h0d02, 16'h0d01, 16'h0d00, 16'h0cff, 16'h0cfe, 16'h0cfd, 16'h0cfc, 16'h0cfb, 16'h0cfa, 16'h0cf9, 16'h0cf8, 16'h0cf7, 16'h0cf6, 16'h0cf5, 16'h0cf4, 16'h0cf3, 16'h0cf2, 16'h0cf1, 16'h0cf0, 16'h0cef, 16'h0cee, 16'h0ced, 16'h0cec, 16'h0ceb, 16'h0cea, 16'h0ce9, 16'h0ce8, 16'h0ce7, 16'h0ce6, 16'h0ce5, 16'h0ce4, 16'h0ce3, 16'h0ce2},
                                {16'h0ce1, 16'h0ce0, 16'h0cdf, 16'h0cde, 16'h0cdd, 16'h0cdc, 16'h0cdb, 16'h0cda, 16'h0cd9, 16'h0cd8, 16'h0cd7, 16'h0cd6, 16'h0cd5, 16'h0cd4, 16'h0cd3, 16'h0cd2, 16'h0cd1, 16'h0cd0, 16'h0ccf, 16'h0cce, 16'h0ccd, 16'h0ccc, 16'h0ccb, 16'h0cca, 16'h0cc9, 16'h0cc8, 16'h0cc7, 16'h0cc6, 16'h0cc5, 16'h0cc4, 16'h0cc3, 16'h0cc2, 16'h0cc1, 16'h0cc0, 16'h0cbf, 16'h0cbe, 16'h0cbd, 16'h0cbc, 16'h0cbb, 16'h0cba, 16'h0cb9, 16'h0cb8, 16'h0cb7, 16'h0cb6, 16'h0cb5, 16'h0cb4, 16'h0cb3, 16'h0cb2, 16'h0cb1, 16'h0cb0, 16'h0caf, 16'h0cae, 16'h0cad, 16'h0cac, 16'h0cab, 16'h0caa, 16'h0ca9, 16'h0ca8, 16'h0ca7, 16'h0ca6, 16'h0ca5, 16'h0ca4, 16'h0ca3, 16'h0ca2},
                                {16'h0ca1, 16'h0ca0, 16'h0c9f, 16'h0c9e, 16'h0c9d, 16'h0c9c, 16'h0c9b, 16'h0c9a, 16'h0c99, 16'h0c98, 16'h0c97, 16'h0c96, 16'h0c95, 16'h0c94, 16'h0c93, 16'h0c92, 16'h0c91, 16'h0c90, 16'h0c8f, 16'h0c8e, 16'h0c8d, 16'h0c8c, 16'h0c8b, 16'h0c8a, 16'h0c89, 16'h0c88, 16'h0c87, 16'h0c86, 16'h0c85, 16'h0c84, 16'h0c83, 16'h0c82, 16'h0c81, 16'h0c80, 16'h0c7f, 16'h0c7e, 16'h0c7d, 16'h0c7c, 16'h0c7b, 16'h0c7a, 16'h0c79, 16'h0c78, 16'h0c77, 16'h0c76, 16'h0c75, 16'h0c74, 16'h0c73, 16'h0c72, 16'h0c71, 16'h0c70, 16'h0c6f, 16'h0c6e, 16'h0c6d, 16'h0c6c, 16'h0c6b, 16'h0c6a, 16'h0c69, 16'h0c68, 16'h0c67, 16'h0c66, 16'h0c65, 16'h0c64, 16'h0c63, 16'h0c62},
                                {16'h0c61, 16'h0c60, 16'h0c5f, 16'h0c5e, 16'h0c5d, 16'h0c5c, 16'h0c5b, 16'h0c5a, 16'h0c59, 16'h0c58, 16'h0c57, 16'h0c56, 16'h0c55, 16'h0c54, 16'h0c53, 16'h0c52, 16'h0c51, 16'h0c50, 16'h0c4f, 16'h0c4e, 16'h0c4d, 16'h0c4c, 16'h0c4b, 16'h0c4a, 16'h0c49, 16'h0c48, 16'h0c47, 16'h0c46, 16'h0c45, 16'h0c44, 16'h0c43, 16'h0c42, 16'h0c41, 16'h0c40, 16'h0c3f, 16'h0c3e, 16'h0c3d, 16'h0c3c, 16'h0c3b, 16'h0c3a, 16'h0c39, 16'h0c38, 16'h0c37, 16'h0c36, 16'h0c35, 16'h0c34, 16'h0c33, 16'h0c32, 16'h0c31, 16'h0c30, 16'h0c2f, 16'h0c2e, 16'h0c2d, 16'h0c2c, 16'h0c2b, 16'h0c2a, 16'h0c29, 16'h0c28, 16'h0c27, 16'h0c26, 16'h0c25, 16'h0c24, 16'h0c23, 16'h0c22},
                                {16'h0c21, 16'h0c20, 16'h0c1f, 16'h0c1e, 16'h0c1d, 16'h0c1c, 16'h0c1b, 16'h0c1a, 16'h0c19, 16'h0c18, 16'h0c17, 16'h0c16, 16'h0c15, 16'h0c14, 16'h0c13, 16'h0c12, 16'h0c11, 16'h0c10, 16'h0c0f, 16'h0c0e, 16'h0c0d, 16'h0c0c, 16'h0c0b, 16'h0c0a, 16'h0c09, 16'h0c08, 16'h0c07, 16'h0c06, 16'h0c05, 16'h0c04, 16'h0c03, 16'h0c02, 16'h0c01, 16'h0c00, 16'h0bff, 16'h0bfe, 16'h0bfd, 16'h0bfc, 16'h0bfb, 16'h0bfa, 16'h0bf9, 16'h0bf8, 16'h0bf7, 16'h0bf6, 16'h0bf5, 16'h0bf4, 16'h0bf3, 16'h0bf2, 16'h0bf1, 16'h0bf0, 16'h0bef, 16'h0bee, 16'h0bed, 16'h0bec, 16'h0beb, 16'h0bea, 16'h0be9, 16'h0be8, 16'h0be7, 16'h0be6, 16'h0be5, 16'h0be4, 16'h0be3, 16'h0be2},
                                {16'h0be1, 16'h0be0, 16'h0bdf, 16'h0bde, 16'h0bdd, 16'h0bdc, 16'h0bdb, 16'h0bda, 16'h0bd9, 16'h0bd8, 16'h0bd7, 16'h0bd6, 16'h0bd5, 16'h0bd4, 16'h0bd3, 16'h0bd2, 16'h0bd1, 16'h0bd0, 16'h0bcf, 16'h0bce, 16'h0bcd, 16'h0bcc, 16'h0bcb, 16'h0bca, 16'h0bc9, 16'h0bc8, 16'h0bc7, 16'h0bc6, 16'h0bc5, 16'h0bc4, 16'h0bc3, 16'h0bc2, 16'h0bc1, 16'h0bc0, 16'h0bbf, 16'h0bbe, 16'h0bbd, 16'h0bbc, 16'h0bbb, 16'h0bba, 16'h0bb9, 16'h0bb8, 16'h0bb7, 16'h0bb6, 16'h0bb5, 16'h0bb4, 16'h0bb3, 16'h0bb2, 16'h0bb1, 16'h0bb0, 16'h0baf, 16'h0bae, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad},
                                {16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad},
                                {16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad},
                                {16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad},
                                {16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad},
                                {16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad},
                                {16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad},
                                {16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad},
                                {16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad},
                                {16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad},
                                {16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad},
                                {16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad},
                                {16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bad, 16'h0bac, 16'h0bab, 16'h0baa, 16'h0ba9, 16'h0ba8},
                                {16'h0ba7, 16'h0ba6, 16'h0ba5, 16'h0ba4, 16'h0ba3, 16'h0ba2, 16'h0ba1, 16'h0ba0, 16'h0b9f, 16'h0b9e, 16'h0b9d, 16'h0b9c, 16'h0b9b, 16'h0b9a, 16'h0b99, 16'h0b98, 16'h0b97, 16'h0b96, 16'h0b95, 16'h0b94, 16'h0b93, 16'h0b92, 16'h0b91, 16'h0b90, 16'h0b8f, 16'h0b8e, 16'h0b8d, 16'h0b8c, 16'h0b8b, 16'h0b8a, 16'h0b89, 16'h0b88, 16'h0b87, 16'h0b86, 16'h0b85, 16'h0b84, 16'h0b83, 16'h0b82, 16'h0b81, 16'h0b80, 16'h0b7f, 16'h0b7e, 16'h0b7d, 16'h0b7c, 16'h0b7b, 16'h0b7a, 16'h0b79, 16'h0b78, 16'h0b77, 16'h0b76, 16'h0b75, 16'h0b74, 16'h0b73, 16'h0b72, 16'h0b71, 16'h0b70, 16'h0b6f, 16'h0b6e, 16'h0b6d, 16'h0b6c, 16'h0b6b, 16'h0b6a, 16'h0b69, 16'h0b68},
                                {16'h0b67, 16'h0b66, 16'h0b65, 16'h0b64, 16'h0b63, 16'h0b62, 16'h0b61, 16'h0b60, 16'h0b5f, 16'h0b5e, 16'h0b5d, 16'h0b5c, 16'h0b5b, 16'h0b5a, 16'h0b59, 16'h0b58, 16'h0b57, 16'h0b56, 16'h0b55, 16'h0b54, 16'h0b53, 16'h0b52, 16'h0b51, 16'h0b50, 16'h0b4f, 16'h0b4e, 16'h0b4d, 16'h0b4c, 16'h0b4b, 16'h0b4a, 16'h0b49, 16'h0b48, 16'h0b47, 16'h0b46, 16'h0b45, 16'h0b44, 16'h0b43, 16'h0b42, 16'h0b41, 16'h0b40, 16'h0b3f, 16'h0b3e, 16'h0b3d, 16'h0b3c, 16'h0b3b, 16'h0b3a, 16'h0b39, 16'h0b38, 16'h0b37, 16'h0b36, 16'h0b35, 16'h0b34, 16'h0b33, 16'h0b32, 16'h0b31, 16'h0b30, 16'h0b2f, 16'h0b2e, 16'h0b2d, 16'h0b2c, 16'h0b2b, 16'h0b2a, 16'h0b29, 16'h0b28},
                                {16'h0b27, 16'h0b26, 16'h0b25, 16'h0b24, 16'h0b23, 16'h0b22, 16'h0b21, 16'h0b20, 16'h0b1f, 16'h0b1e, 16'h0b1d, 16'h0b1c, 16'h0b1b, 16'h0b1a, 16'h0b19, 16'h0b18, 16'h0b17, 16'h0b16, 16'h0b15, 16'h0b14, 16'h0b13, 16'h0b12, 16'h0b11, 16'h0b10, 16'h0b0f, 16'h0b0e, 16'h0b0d, 16'h0b0c, 16'h0b0b, 16'h0b0a, 16'h0b09, 16'h0b08, 16'h0b07, 16'h0b06, 16'h0b05, 16'h0b04, 16'h0b03, 16'h0b02, 16'h0b01, 16'h0b00, 16'h0aff, 16'h0afe, 16'h0afd, 16'h0afc, 16'h0afb, 16'h0afa, 16'h0af9, 16'h0af8, 16'h0af7, 16'h0af6, 16'h0af5, 16'h0af4, 16'h0af3, 16'h0af2, 16'h0af1, 16'h0af0, 16'h0aef, 16'h0aee, 16'h0aed, 16'h0aec, 16'h0aeb, 16'h0aea, 16'h0ae9, 16'h0ae8},
                                {16'h0ae7, 16'h0ae6, 16'h0ae5, 16'h0ae4, 16'h0ae3, 16'h0ae2, 16'h0ae1, 16'h0ae0, 16'h0adf, 16'h0ade, 16'h0add, 16'h0adc, 16'h0adb, 16'h0ada, 16'h0ad9, 16'h0ad8, 16'h0ad7, 16'h0ad6, 16'h0ad5, 16'h0ad4, 16'h0ad3, 16'h0ad2, 16'h0ad1, 16'h0ad0, 16'h0acf, 16'h0ace, 16'h0acd, 16'h0acc, 16'h0acb, 16'h0aca, 16'h0ac9, 16'h0ac8, 16'h0ac7, 16'h0ac6, 16'h0ac5, 16'h0ac4, 16'h0ac3, 16'h0ac2, 16'h0ac1, 16'h0ac0, 16'h0abf, 16'h0abe, 16'h0abd, 16'h0abc, 16'h0abb, 16'h0aba, 16'h0ab9, 16'h0ab8, 16'h0ab7, 16'h0ab6, 16'h0ab5, 16'h0ab4, 16'h0ab3, 16'h0ab2, 16'h0ab1, 16'h0ab0, 16'h0aaf, 16'h0aae, 16'h0aad, 16'h0aac, 16'h0aab, 16'h0aaa, 16'h0aa9, 16'h0aa8},
                                {16'h0aa7, 16'h0aa6, 16'h0aa5, 16'h0aa4, 16'h0aa3, 16'h0aa2, 16'h0aa1, 16'h0aa0, 16'h0a9f, 16'h0a9e, 16'h0a9d, 16'h0a9c, 16'h0a9b, 16'h0a9a, 16'h0a99, 16'h0a98, 16'h0a97, 16'h0a96, 16'h0a95, 16'h0a94, 16'h0a93, 16'h0a92, 16'h0a91, 16'h0a90, 16'h0a8f, 16'h0a8e, 16'h0a8d, 16'h0a8c, 16'h0a8b, 16'h0a8a, 16'h0a89, 16'h0a88, 16'h0a87, 16'h0a86, 16'h0a85, 16'h0a84, 16'h0a83, 16'h0a82, 16'h0a81, 16'h0a80, 16'h0a7f, 16'h0a7e, 16'h0a7d, 16'h0a7c, 16'h0a7b, 16'h0a7a, 16'h0a79, 16'h0a78, 16'h0a77, 16'h0a76, 16'h0a75, 16'h0a74, 16'h0a73, 16'h0a72, 16'h0a71, 16'h0a70, 16'h0a6f, 16'h0a6e, 16'h0a6d, 16'h0a6c, 16'h0a6b, 16'h0a6a, 16'h0a69, 16'h0a68},
                                {16'h0a67, 16'h0a66, 16'h0a65, 16'h0a64, 16'h0a63, 16'h0a62, 16'h0a61, 16'h0a60, 16'h0a5f, 16'h0a5e, 16'h0a5d, 16'h0a5c, 16'h0a5b, 16'h0a5a, 16'h0a59, 16'h0a58, 16'h0a57, 16'h0a56, 16'h0a55, 16'h0a54, 16'h0a53, 16'h0a52, 16'h0a51, 16'h0a50, 16'h0a4f, 16'h0a4e, 16'h0a4d, 16'h0a4c, 16'h0a4b, 16'h0a4a, 16'h0a49, 16'h0a48, 16'h0a47, 16'h0a46, 16'h0a45, 16'h0a44, 16'h0a43, 16'h0a42, 16'h0a41, 16'h0a40, 16'h0a3f, 16'h0a3e, 16'h0a3d, 16'h0a3c, 16'h0a3b, 16'h0a3a, 16'h0a39, 16'h0a38, 16'h0a37, 16'h0a36, 16'h0a35, 16'h0a34, 16'h0a33, 16'h0a32, 16'h0a31, 16'h0a30, 16'h0a2f, 16'h0a2e, 16'h0a2d, 16'h0a2c, 16'h0a2b, 16'h0a2a, 16'h0a29, 16'h0a28},
                                {16'h0a27, 16'h0a26, 16'h0a25, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24},
                                {16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24},
                                {16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24},
                                {16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24},
                                {16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24},
                                {16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24},
                                {16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24},
                                {16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24},
                                {16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24},
                                {16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24},
                                {16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24},
                                {16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24},
                                {16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a24, 16'h0a23, 16'h0a22, 16'h0a21, 16'h0a20, 16'h0a1f, 16'h0a1e, 16'h0a1d, 16'h0a1c, 16'h0a1b, 16'h0a1a, 16'h0a19, 16'h0a18, 16'h0a17, 16'h0a16, 16'h0a15, 16'h0a14, 16'h0a13, 16'h0a12, 16'h0a11, 16'h0a10, 16'h0a0f, 16'h0a0e, 16'h0a0d, 16'h0a0c, 16'h0a0b, 16'h0a0a, 16'h0a09, 16'h0a08, 16'h0a07, 16'h0a06, 16'h0a05, 16'h0a04, 16'h0a03, 16'h0a02, 16'h0a01, 16'h0a00, 16'h09ff, 16'h09fe, 16'h09fd, 16'h09fc, 16'h09fb, 16'h09fa, 16'h09f9, 16'h09f8, 16'h09f7, 16'h09f6, 16'h09f5, 16'h09f4, 16'h09f3, 16'h09f2, 16'h09f1, 16'h09f0, 16'h09ef, 16'h09ee, 16'h09ed},
                                {16'h09ec, 16'h09eb, 16'h09ea, 16'h09e9, 16'h09e8, 16'h09e7, 16'h09e6, 16'h09e5, 16'h09e4, 16'h09e3, 16'h09e2, 16'h09e1, 16'h09e0, 16'h09df, 16'h09de, 16'h09dd, 16'h09dc, 16'h09db, 16'h09da, 16'h09d9, 16'h09d8, 16'h09d7, 16'h09d6, 16'h09d5, 16'h09d4, 16'h09d3, 16'h09d2, 16'h09d1, 16'h09d0, 16'h09cf, 16'h09ce, 16'h09cd, 16'h09cc, 16'h09cb, 16'h09ca, 16'h09c9, 16'h09c8, 16'h09c7, 16'h09c6, 16'h09c5, 16'h09c4, 16'h09c3, 16'h09c2, 16'h09c1, 16'h09c0, 16'h09bf, 16'h09be, 16'h09bd, 16'h09bc, 16'h09bb, 16'h09ba, 16'h09b9, 16'h09b8, 16'h09b7, 16'h09b6, 16'h09b5, 16'h09b4, 16'h09b3, 16'h09b2, 16'h09b1, 16'h09b0, 16'h09af, 16'h09ae, 16'h09ad},
                                {16'h09ac, 16'h09ab, 16'h09aa, 16'h09a9, 16'h09a8, 16'h09a7, 16'h09a6, 16'h09a5, 16'h09a4, 16'h09a3, 16'h09a2, 16'h09a1, 16'h09a0, 16'h099f, 16'h099e, 16'h099d, 16'h099c, 16'h099b, 16'h099a, 16'h0999, 16'h0998, 16'h0997, 16'h0996, 16'h0995, 16'h0994, 16'h0993, 16'h0992, 16'h0991, 16'h0990, 16'h098f, 16'h098e, 16'h098d, 16'h098c, 16'h098b, 16'h098a, 16'h0989, 16'h0988, 16'h0987, 16'h0986, 16'h0985, 16'h0984, 16'h0983, 16'h0982, 16'h0981, 16'h0980, 16'h097f, 16'h097e, 16'h097d, 16'h097c, 16'h097b, 16'h097a, 16'h0979, 16'h0978, 16'h0977, 16'h0976, 16'h0975, 16'h0974, 16'h0973, 16'h0972, 16'h0971, 16'h0970, 16'h096f, 16'h096e, 16'h096d},
                                {16'h096c, 16'h096b, 16'h096a, 16'h0969, 16'h0968, 16'h0967, 16'h0966, 16'h0965, 16'h0964, 16'h0963, 16'h0962, 16'h0961, 16'h0960, 16'h095f, 16'h095e, 16'h095d, 16'h095c, 16'h095b, 16'h095a, 16'h0959, 16'h0958, 16'h0957, 16'h0956, 16'h0955, 16'h0954, 16'h0953, 16'h0952, 16'h0951, 16'h0950, 16'h094f, 16'h094e, 16'h094d, 16'h094c, 16'h094b, 16'h094a, 16'h0949, 16'h0948, 16'h0947, 16'h0946, 16'h0945, 16'h0944, 16'h0943, 16'h0942, 16'h0941, 16'h0940, 16'h093f, 16'h093e, 16'h093d, 16'h093c, 16'h093b, 16'h093a, 16'h0939, 16'h0938, 16'h0937, 16'h0936, 16'h0935, 16'h0934, 16'h0933, 16'h0932, 16'h0931, 16'h0930, 16'h092f, 16'h092e, 16'h092d},
                                {16'h092c, 16'h092b, 16'h092a, 16'h0929, 16'h0928, 16'h0927, 16'h0926, 16'h0925, 16'h0924, 16'h0923, 16'h0922, 16'h0921, 16'h0920, 16'h091f, 16'h091e, 16'h091d, 16'h091c, 16'h091b, 16'h091a, 16'h0919, 16'h0918, 16'h0917, 16'h0916, 16'h0915, 16'h0914, 16'h0913, 16'h0912, 16'h0911, 16'h0910, 16'h090f, 16'h090e, 16'h090d, 16'h090c, 16'h090b, 16'h090a, 16'h0909, 16'h0908, 16'h0907, 16'h0906, 16'h0905, 16'h0904, 16'h0903, 16'h0902, 16'h0901, 16'h0900, 16'h08ff, 16'h08fe, 16'h08fd, 16'h08fc, 16'h08fb, 16'h08fa, 16'h08f9, 16'h08f8, 16'h08f7, 16'h08f6, 16'h08f5, 16'h08f4, 16'h08f3, 16'h08f2, 16'h08f1, 16'h08f0, 16'h08ef, 16'h08ee, 16'h08ed},
                                {16'h08ec, 16'h08eb, 16'h08ea, 16'h08e9, 16'h08e8, 16'h08e7, 16'h08e6, 16'h08e5, 16'h08e4, 16'h08e3, 16'h08e2, 16'h08e1, 16'h08e0, 16'h08df, 16'h08de, 16'h08dd, 16'h08dc, 16'h08db, 16'h08da, 16'h08d9, 16'h08d8, 16'h08d7, 16'h08d6, 16'h08d5, 16'h08d4, 16'h08d3, 16'h08d2, 16'h08d1, 16'h08d0, 16'h08cf, 16'h08ce, 16'h08cd, 16'h08cc, 16'h08cb, 16'h08ca, 16'h08c9, 16'h08c8, 16'h08c7, 16'h08c6, 16'h08c5, 16'h08c4, 16'h08c3, 16'h08c2, 16'h08c1, 16'h08c0, 16'h08bf, 16'h08be, 16'h08bd, 16'h08bc, 16'h08bb, 16'h08ba, 16'h08b9, 16'h08b8, 16'h08b7, 16'h08b6, 16'h08b5, 16'h08b4, 16'h08b3, 16'h08b2, 16'h08b1, 16'h08b0, 16'h08af, 16'h08ae, 16'h0a10},
                                {16'h0a11, 16'h0a12, 16'h0a13, 16'h0a14, 16'h0a15, 16'h0a16, 16'h0a17, 16'h0a18, 16'h0a19, 16'h0a1a, 16'h0a1b, 16'h0a1c, 16'h0a1d, 16'h0a1e, 16'h0a1f, 16'h0a20, 16'h0a21, 16'h0a22, 16'h0a23, 16'h0a24, 16'h0a25, 16'h0a26, 16'h0a27, 16'h0a28, 16'h0a29, 16'h0a2a, 16'h0a2b, 16'h0a2c, 16'h0a2d, 16'h0a2e, 16'h0a2f, 16'h0a30, 16'h0a31, 16'h0a32, 16'h0a33, 16'h0a34, 16'h0a35, 16'h0a36, 16'h0a37, 16'h0a38, 16'h0a39, 16'h0a3a, 16'h0a3b, 16'h0a3c, 16'h0a3d, 16'h0a3e, 16'h0a3f, 16'h0a40, 16'h0a41, 16'h0a42, 16'h0a43, 16'h0a44, 16'h0a45, 16'h0a46, 16'h0a47, 16'h0a48, 16'h0a49, 16'h0a4a, 16'h0a4b, 16'h0a4c, 16'h0a4d, 16'h0a4e, 16'h0a4f, 16'h0a50},
                                {16'h0a51, 16'h0a52, 16'h0a53, 16'h0a54, 16'h0a55, 16'h0a56, 16'h0a57, 16'h0a58, 16'h0a59, 16'h0a5a, 16'h0a5b, 16'h0a5c, 16'h0a5d, 16'h0a5e, 16'h0a5f, 16'h0a60, 16'h0a61, 16'h0a62, 16'h0a63, 16'h0a64, 16'h0a65, 16'h0a66, 16'h0a67, 16'h0a68, 16'h0a69, 16'h0a6a, 16'h0a6b, 16'h0a6c, 16'h0a6d, 16'h0a6e, 16'h0a6f, 16'h0a70, 16'h0a71, 16'h0a72, 16'h0a73, 16'h0a74, 16'h0a75, 16'h0a76, 16'h0a77, 16'h0a78, 16'h0a79, 16'h0a7a, 16'h0a7b, 16'h0a7c, 16'h0a7d, 16'h0a7e, 16'h0a7f, 16'h0a80, 16'h0a81, 16'h0a82, 16'h0a83, 16'h0a84, 16'h0a85, 16'h0a86, 16'h0a87, 16'h0a88, 16'h0a89, 16'h0a8a, 16'h0a8b, 16'h0a8c, 16'h0a8d, 16'h0a8e, 16'h0a8f, 16'h0a90},
                                {16'h0a91, 16'h0a92, 16'h0a93, 16'h0a94, 16'h0a95, 16'h0a96, 16'h0a97, 16'h0a98, 16'h0a99, 16'h0a9a, 16'h0a9b, 16'h0a9c, 16'h0a9d, 16'h0a9e, 16'h0a9f, 16'h0aa0, 16'h0aa1, 16'h0aa2, 16'h0aa3, 16'h0aa4, 16'h0aa5, 16'h0aa6, 16'h0aa7, 16'h0aa8, 16'h0aa9, 16'h0aaa, 16'h0aab, 16'h0aac, 16'h0aad, 16'h0aae, 16'h0aaf, 16'h0ab0, 16'h0ab1, 16'h0ab2, 16'h0ab3, 16'h0ab4, 16'h0ab5, 16'h0ab6, 16'h0ab7, 16'h0ab8, 16'h0ab9, 16'h0aba, 16'h0abb, 16'h0abc, 16'h0abd, 16'h0abe, 16'h0abf, 16'h0ac0, 16'h0ac1, 16'h0ac2, 16'h0ac3, 16'h0ac4, 16'h0ac5, 16'h0ac6, 16'h0ac7, 16'h0ac8, 16'h0ac9, 16'h0aca, 16'h0acb, 16'h0acc, 16'h0acd, 16'h0ace, 16'h0acf, 16'h0ad0},
                                {16'h0ad1, 16'h0ad2, 16'h0ad3, 16'h0ad4, 16'h0ad5, 16'h0ad6, 16'h0ad7, 16'h0ad8, 16'h0ad9, 16'h0ada, 16'h0adb, 16'h0adc, 16'h0add, 16'h0ade, 16'h0adf, 16'h0ae0, 16'h0ae1, 16'h0ae2, 16'h0ae3, 16'h0ae4, 16'h0ae5, 16'h0ae6, 16'h0ae7, 16'h0ae8, 16'h0ae9, 16'h0aea, 16'h0aeb, 16'h0aec, 16'h0aed, 16'h0aee, 16'h0aef, 16'h0af0, 16'h0af1, 16'h0af2, 16'h0af3, 16'h0af4, 16'h0af5, 16'h0af6, 16'h0af7, 16'h0af8, 16'h0af9, 16'h0afa, 16'h0afb, 16'h0afc, 16'h0afd, 16'h0afe, 16'h0aff, 16'h0b00, 16'h0b01, 16'h0b02, 16'h0b03, 16'h0b04, 16'h0b05, 16'h0b06, 16'h0b07, 16'h0b08, 16'h0b09, 16'h0b0a, 16'h0b0b, 16'h0b0c, 16'h0b0d, 16'h0b0e, 16'h0b0f, 16'h0b10},
                                {16'h0b11, 16'h0b12, 16'h0b13, 16'h0b14, 16'h0b15, 16'h0b16, 16'h0b17, 16'h0b18, 16'h0b19, 16'h0b1a, 16'h0b1b, 16'h0b1c, 16'h0b1d, 16'h0b1e, 16'h0b1f, 16'h0b20, 16'h0b21, 16'h0b22, 16'h0b23, 16'h0b24, 16'h0b25, 16'h0b26, 16'h0b27, 16'h0b28, 16'h0b29, 16'h0b2a, 16'h0b2b, 16'h0b2c, 16'h0b2d, 16'h0b2e, 16'h0b2f, 16'h0b30, 16'h0b31, 16'h0b32, 16'h0b33, 16'h0b34, 16'h0b35, 16'h0b36, 16'h0b37, 16'h0b38, 16'h0b39, 16'h0b3a, 16'h0b3b, 16'h0b3c, 16'h0b3d, 16'h0b3e, 16'h0b3f, 16'h0b40, 16'h0b41, 16'h0b42, 16'h0b43, 16'h0b44, 16'h0b45, 16'h0b46, 16'h0b47, 16'h0b48, 16'h0b49, 16'h0b4a, 16'h0b4b, 16'h0b4c, 16'h0b4d, 16'h0b4e, 16'h0b4f, 16'h0b50},
                                {16'h0b51, 16'h0b52, 16'h0b53, 16'h0b54, 16'h0b55, 16'h0b56, 16'h0b57, 16'h0b58, 16'h0b59, 16'h0b5a, 16'h0b5b, 16'h0b5c, 16'h0b5d, 16'h0b5e, 16'h0b5f, 16'h0b60, 16'h0b61, 16'h0b62, 16'h0b63, 16'h0b64, 16'h0b65, 16'h0b66, 16'h0b67, 16'h0b68, 16'h0b69, 16'h0b6a, 16'h0b6b, 16'h0b6c, 16'h0b6d, 16'h0b6e, 16'h0b6f, 16'h0b70, 16'h0b71, 16'h0b72, 16'h0b73, 16'h0b74, 16'h0b75, 16'h0b76, 16'h0b77, 16'h0b78, 16'h0b79, 16'h0b7a, 16'h0b7b, 16'h0b7c, 16'h0b7d, 16'h0b7e, 16'h0b7f, 16'h0b80, 16'h0b81, 16'h0b82, 16'h0b83, 16'h0b84, 16'h0b85, 16'h0b86, 16'h0b87, 16'h0b88, 16'h0b89, 16'h0b8a, 16'h0b8b, 16'h0b8c, 16'h0b8d, 16'h0b8e, 16'h0b8f, 16'h0b90},
                                {16'h0b91, 16'h0b92, 16'h0b93, 16'h0b94, 16'h0b95, 16'h0b96, 16'h0b97, 16'h0b98, 16'h0b99, 16'h0b9a, 16'h0b9b, 16'h0b9c, 16'h0b9d, 16'h0b9e, 16'h0b9f, 16'h0ba0, 16'h0ba1, 16'h0ba2, 16'h0ba3, 16'h0ba4, 16'h0ba5, 16'h0ba6, 16'h0ba7, 16'h0ba8, 16'h0ba9, 16'h0baa, 16'h0bab, 16'h0bac, 16'h0bad, 16'h0bae, 16'h0baf, 16'h0bb0, 16'h0bb1, 16'h0bb2, 16'h0bb3, 16'h0bb4, 16'h0bb5, 16'h0bb6, 16'h0bb7, 16'h0bb8, 16'h0bb9, 16'h0bba, 16'h0bbb, 16'h0bbc, 16'h0bbd, 16'h0bbe, 16'h0bbf, 16'h0bc0, 16'h0bc1, 16'h0bc2, 16'h0bc3, 16'h0bc4, 16'h0bc5, 16'h0bc6, 16'h0bc7, 16'h0bc8, 16'h0bc9, 16'h0bca, 16'h0bcb, 16'h0bcc, 16'h0bcd, 16'h0bce, 16'h0bcf, 16'h0bd0},
                                {16'h0bd1, 16'h0bd2, 16'h0bd3, 16'h0bd4, 16'h0bd5, 16'h0bd6, 16'h0bd7, 16'h0bd8, 16'h0bd9, 16'h0bda, 16'h0bdb, 16'h0bdc, 16'h0bdd, 16'h0bde, 16'h0bdf, 16'h0be0, 16'h0be1, 16'h0be2, 16'h0be3, 16'h0be4, 16'h0be5, 16'h0be6, 16'h0be7, 16'h0be8, 16'h0be9, 16'h0bea, 16'h0beb, 16'h0bec, 16'h0bed, 16'h0bee, 16'h0bef, 16'h0bf0, 16'h0bf1, 16'h0bf2, 16'h0bf3, 16'h0bf4, 16'h0bf5, 16'h0bf6, 16'h0bf7, 16'h0bf8, 16'h0bf9, 16'h0bfa, 16'h0bfb, 16'h0bfc, 16'h0bfd, 16'h0bfe, 16'h0bff, 16'h0c00, 16'h0c01, 16'h0c02, 16'h0c03, 16'h0c04, 16'h0c05, 16'h0c06, 16'h0c07, 16'h0c08, 16'h0c09, 16'h0c0a, 16'h0c0b, 16'h0c0c, 16'h0c0d, 16'h0c0e, 16'h0c0f, 16'h0c10},
                                {16'h0c11, 16'h0c12, 16'h0c13, 16'h0c14, 16'h0c15, 16'h0c16, 16'h0c17, 16'h0c18, 16'h0c19, 16'h0c1a, 16'h0c1b, 16'h0c1c, 16'h0c1d, 16'h0c1e, 16'h0c1f, 16'h0c20, 16'h0c21, 16'h0c22, 16'h0c23, 16'h0c24, 16'h0c25, 16'h0c26, 16'h0c27, 16'h0c28, 16'h0c29, 16'h0c2a, 16'h0c2b, 16'h0c2c, 16'h0c2d, 16'h0c2e, 16'h0c2f, 16'h0c30, 16'h0c31, 16'h0c32, 16'h0c33, 16'h0c34, 16'h0c35, 16'h0c36, 16'h0c37, 16'h0c38, 16'h0c39, 16'h0c3a, 16'h0c3b, 16'h0c3c, 16'h0c3d, 16'h0c3e, 16'h0c3f, 16'h0c40, 16'h0c41, 16'h0c42, 16'h0c43, 16'h0c44, 16'h0c45, 16'h0c46, 16'h0c47, 16'h0c48, 16'h0c49, 16'h0c4a, 16'h0c4b, 16'h0c4c, 16'h0c4d, 16'h0c4e, 16'h0c4f, 16'h0c50},
                                {16'h0c51, 16'h0c52, 16'h0c53, 16'h0c54, 16'h0c55, 16'h0c56, 16'h0c57, 16'h0c58, 16'h0c59, 16'h0c5a, 16'h0c5b, 16'h0c5c, 16'h0c5d, 16'h0c5e, 16'h0c5f, 16'h0c60, 16'h0c61, 16'h0c62, 16'h0c63, 16'h0c64, 16'h0c65, 16'h0c66, 16'h0c67, 16'h0c68, 16'h0c69, 16'h0c6a, 16'h0c6b, 16'h0c6c, 16'h0c6d, 16'h0c6e, 16'h0c6f, 16'h0c70, 16'h0c71, 16'h0c72, 16'h0c73, 16'h0c74, 16'h0c75, 16'h0c76, 16'h0c77, 16'h0c78, 16'h0c79, 16'h0c7a, 16'h0c7b, 16'h0c7c, 16'h0c7d, 16'h0c7e, 16'h0c7f, 16'h0c80, 16'h0c81, 16'h0c82, 16'h0c83, 16'h0c84, 16'h0c85, 16'h0c86, 16'h0c87, 16'h0c88, 16'h0c89, 16'h0c8a, 16'h0c8b, 16'h0c8c, 16'h0c8d, 16'h0c8e, 16'h0c8f, 16'h0c90},
                                {16'h0c91, 16'h0c92, 16'h0c93, 16'h0c94, 16'h0c95, 16'h0c96, 16'h0c97, 16'h0c98, 16'h0c99, 16'h0c9a, 16'h0c9b, 16'h0c9c, 16'h0c9d, 16'h0c9e, 16'h0c9f, 16'h0ca0, 16'h0ca1, 16'h0ca2, 16'h0ca3, 16'h0ca4, 16'h0ca5, 16'h0ca6, 16'h0ca7, 16'h0ca8, 16'h0ca9, 16'h0caa, 16'h0cab, 16'h0cac, 16'h0cad, 16'h0cae, 16'h0caf, 16'h0cb0, 16'h0cb1, 16'h0cb2, 16'h0cb3, 16'h0cb4, 16'h0cb5, 16'h0cb6, 16'h0cb7, 16'h0cb8, 16'h0cb9, 16'h0cba, 16'h0cbb, 16'h0cbc, 16'h0cbd, 16'h0cbe, 16'h0cbf, 16'h0cc0, 16'h0cc1, 16'h0cc2, 16'h0cc3, 16'h0cc4, 16'h0cc5, 16'h0cc6, 16'h0cc7, 16'h0cc8, 16'h0cc9, 16'h0cca, 16'h0ccb, 16'h0ccc, 16'h0ccd, 16'h0cce, 16'h0ccf, 16'h0cd0},
                                {16'h0cd1, 16'h0cd2, 16'h0cd3, 16'h0cd4, 16'h0cd5, 16'h0cd6, 16'h0cd7, 16'h0cd8, 16'h0cd9, 16'h0cda, 16'h0cdb, 16'h0cdc, 16'h0cdd, 16'h0cde, 16'h0cdf, 16'h0ce0, 16'h0ce1, 16'h0ce2, 16'h0ce3, 16'h0ce4, 16'h0ce5, 16'h0ce6, 16'h0ce7, 16'h0ce8, 16'h0ce9, 16'h0cea, 16'h0ceb, 16'h0cec, 16'h0ced, 16'h0cee, 16'h0cef, 16'h0cf0, 16'h0cf1, 16'h0cf2, 16'h0cf3, 16'h0cf4, 16'h0cf5, 16'h0cf6, 16'h0cf7, 16'h0cf8, 16'h0cf9, 16'h0cfa, 16'h0cfb, 16'h0cfc, 16'h0cfd, 16'h0cfe, 16'h0cff, 16'h0d00, 16'h0d01, 16'h0d02, 16'h0d03, 16'h0d04, 16'h0d05, 16'h0d06, 16'h0d07, 16'h0d08, 16'h0d09, 16'h0d0a, 16'h0d0b, 16'h0d0c, 16'h0d0d, 16'h0d0e, 16'h0d0f, 16'h0d10},
                                {16'h0d11, 16'h0d12, 16'h0d13, 16'h0d14, 16'h0d15, 16'h0d16, 16'h0d17, 16'h0d18, 16'h0d19, 16'h0d1a, 16'h0d1b, 16'h0d1c, 16'h0d1d, 16'h0d1e, 16'h0d1f, 16'h0d20, 16'h0d21, 16'h0d22, 16'h0d23, 16'h0d24, 16'h0d25, 16'h0d26, 16'h0d27, 16'h0d28, 16'h0d29, 16'h0d2a, 16'h0d2b, 16'h0d2c, 16'h0d2d, 16'h0d2e, 16'h0d2f, 16'h0d30, 16'h0d31, 16'h0d32, 16'h0d33, 16'h0d34, 16'h0d35, 16'h0d36, 16'h0d37, 16'h0d38, 16'h0d39, 16'h0d3a, 16'h0d3b, 16'h0d3c, 16'h0d3d, 16'h0d3e, 16'h0d3f, 16'h0d40, 16'h0d41, 16'h0d42, 16'h0d43, 16'h0d44, 16'h0d45, 16'h0d46, 16'h0d47, 16'h0d48, 16'h0d49, 16'h0d4a, 16'h0d4b, 16'h0d4c, 16'h0d4d, 16'h0d4e, 16'h0d4f, 16'h0d50},
                                {16'h0d51, 16'h0d52, 16'h0d53, 16'h0d54, 16'h0d55, 16'h0d56, 16'h0d57, 16'h0d58, 16'h0d59, 16'h0d5a, 16'h0d5b, 16'h0d5c, 16'h0d5d, 16'h0d5e, 16'h0d7d, 16'h0d81, 16'h0d85, 16'h0d89, 16'h0d8d, 16'h0d91, 16'h0d95, 16'h0d99, 16'h0d9d, 16'h0da1, 16'h0da5, 16'h0da9, 16'h0dad, 16'h0db1, 16'h0db5, 16'h0db9, 16'h0dbd, 16'h0dc1, 16'h0dc5, 16'h0dc9, 16'h0dcd, 16'h0dd1, 16'h0dd5, 16'h0dd9, 16'h0ddd, 16'h0de1, 16'h0de5, 16'h0de9, 16'h0ded, 16'h0df1, 16'h0df5, 16'h0df9, 16'h0dfd, 16'h0e01, 16'h0e05, 16'h0e09, 16'h0e0d, 16'h0e11, 16'h0e15, 16'h0e19, 16'h0e1d, 16'h0e21, 16'h0e25, 16'h0e29, 16'h0e2d, 16'h0e31, 16'h0e35, 16'h0e39, 16'h0e3d, 16'h0e41},
                                {16'h0e45, 16'h0e49, 16'h0e4d, 16'h0e51, 16'h0e55, 16'h0e59, 16'h0e5d, 16'h0e61, 16'h0e65, 16'h0e69, 16'h0e6d, 16'h0e71, 16'h0e75, 16'h0e79, 16'h0e7d, 16'h0e81, 16'h0e85, 16'h0e89, 16'h0e8d, 16'h0e91, 16'h0e95, 16'h0e99, 16'h0e9d, 16'h0ea1, 16'h0ea5, 16'h0ea9, 16'h0ead, 16'h0eb1, 16'h0eb5, 16'h0eb9, 16'h0ebd, 16'h0ec1, 16'h0ec5, 16'h0ec9, 16'h0ecd, 16'h0ed1, 16'h0ed5, 16'h0ed9, 16'h0edd, 16'h0ee1, 16'h0ee5, 16'h0ee9, 16'h0eed, 16'h0ef1, 16'h0ef5, 16'h0ef9, 16'h0efd, 16'h0f01, 16'h0f05, 16'h0f09, 16'h0f0d, 16'h0f11, 16'h0f15, 16'h0f19, 16'h0f1d, 16'h0f21, 16'h0f25, 16'h0f29, 16'h0f2d, 16'h0f31, 16'h0f35, 16'h0f39, 16'h0f3d, 16'h0f41},
                                {16'h0f45, 16'h0f49, 16'h0f4d, 16'h0f51, 16'h0f55, 16'h0f59, 16'h0f5d, 16'h0f61, 16'h0f65, 16'h0f69, 16'h0f6d, 16'h0f71, 16'h0f75, 16'h0f79, 16'h0f7d, 16'h0f81, 16'h0f85, 16'h0f89, 16'h0f8d, 16'h0f91, 16'h0f95, 16'h0f99, 16'h0f9d, 16'h0fa1, 16'h0fa5, 16'h0fa9, 16'h0fad, 16'h0fb1, 16'h0fb5, 16'h0fb9, 16'h0fbd, 16'h0fc1, 16'h0fc5, 16'h0fc9, 16'h0fcd, 16'h0fd1, 16'h0fd5, 16'h0fd9, 16'h0fdd, 16'h0fe1, 16'h0fe5, 16'h0fe9, 16'h0fed, 16'h0ff1, 16'h0ff5, 16'h0ff9, 16'h0ffd, 16'h1001, 16'h1005, 16'h1009, 16'h100d, 16'h1011, 16'h1015, 16'h1019, 16'h101d, 16'h1021, 16'h1025, 16'h1029, 16'h102d, 16'h1031, 16'h1035, 16'h1039, 16'h103d, 16'h1041},
                                {16'h1045, 16'h1049, 16'h104d, 16'h1051, 16'h1055, 16'h1059, 16'h105d, 16'h1061, 16'h1065, 16'h1069, 16'h106d, 16'h1071, 16'h1075, 16'h1079, 16'h107d, 16'h1081, 16'h1085, 16'h1089, 16'h108d, 16'h1091, 16'h1095, 16'h1099, 16'h109d, 16'h10a1, 16'h10a5, 16'h10a9, 16'h10ad, 16'h10b1, 16'h10b5, 16'h10b9, 16'h10bd, 16'h10c1, 16'h10c5, 16'h10c9, 16'h10cd, 16'h10d1, 16'h10d5, 16'h10d9, 16'h10dd, 16'h10e1, 16'h10e5, 16'h10e9, 16'h10ed, 16'h10f1, 16'h10f5, 16'h10f9, 16'h10fd, 16'h1101, 16'h1105, 16'h1109, 16'h110d, 16'h1111, 16'h1115, 16'h1119, 16'h111d, 16'h1121, 16'h1125, 16'h1129, 16'h112d, 16'h1131, 16'h1135, 16'h1139, 16'h113d, 16'h1141},
                                {16'h1145, 16'h1149, 16'h114d, 16'h1151, 16'h1155, 16'h1159, 16'h115d, 16'h1161, 16'h1165, 16'h1169, 16'h116d, 16'h1171, 16'h1175, 16'h1179, 16'h117d, 16'h1181, 16'h1185, 16'h1189, 16'h118d, 16'h1191, 16'h1195, 16'h1199, 16'h119d, 16'h11a1, 16'h11a5, 16'h11a9, 16'h11ad, 16'h11b1, 16'h11b5, 16'h11b9, 16'h11bd, 16'h11c1, 16'h11c5, 16'h11c9, 16'h11cd, 16'h11d1, 16'h11d5, 16'h11d9, 16'h11dd, 16'h11e1, 16'h11e5, 16'h11e9, 16'h11ed, 16'h11f1, 16'h11f5, 16'h11f9, 16'h11fd, 16'h1201, 16'h1205, 16'h1209, 16'h120d, 16'h1211, 16'h1215, 16'h1219, 16'h121d, 16'h1221, 16'h1225, 16'h1229, 16'h122d, 16'h1231, 16'h1235, 16'h1239, 16'h123d, 16'h1241},
                                {16'h1245, 16'h1249, 16'h124d, 16'h1251, 16'h1255, 16'h1259, 16'h125d, 16'h1261, 16'h1265, 16'h1269, 16'h126d, 16'h1271, 16'h1275, 16'h1279, 16'h127d, 16'h1281, 16'h1285, 16'h1289, 16'h128d, 16'h1291, 16'h1295, 16'h1299, 16'h129d, 16'h12a1, 16'h12a5, 16'h12a9, 16'h12ad, 16'h12b1, 16'h12b5, 16'h12b9, 16'h12bd, 16'h12c1, 16'h12c5, 16'h12c9, 16'h12cd, 16'h12d1, 16'h12d5, 16'h12d9, 16'h12dd, 16'h12e1, 16'h12e5, 16'h12e9, 16'h12ed, 16'h12f1, 16'h12f5, 16'h12f9, 16'h12fd, 16'h1301, 16'h1305, 16'h1309, 16'h130d, 16'h1311, 16'h1315, 16'h1319, 16'h131d, 16'h1321, 16'h1325, 16'h1329, 16'h132d, 16'h1331, 16'h1335, 16'h1339, 16'h133d, 16'h1341},
                                {16'h1345, 16'h1349, 16'h134d, 16'h1351, 16'h1355, 16'h1359, 16'h135d, 16'h1361, 16'h1365, 16'h1369, 16'h136d, 16'h1371, 16'h1375, 16'h1379, 16'h137d, 16'h1381, 16'h1385, 16'h1389, 16'h138d, 16'h1391, 16'h1395, 16'h1399, 16'h139d, 16'h13a1, 16'h13a5, 16'h13a9, 16'h13ad, 16'h13b1, 16'h13b5, 16'h13b9, 16'h13bd, 16'h13c1, 16'h13c5, 16'h13c9, 16'h13cd, 16'h13d1, 16'h13d5, 16'h13d9, 16'h13dd, 16'h13e1, 16'h13e5, 16'h13e9, 16'h13ed, 16'h13f1, 16'h13f5, 16'h13f9, 16'h13fd, 16'h1401, 16'h1405, 16'h1409, 16'h140d, 16'h1411, 16'h1415, 16'h1419, 16'h141d, 16'h1421, 16'h1425, 16'h1429, 16'h142d, 16'h1431, 16'h1435, 16'h1439, 16'h143d, 16'h1441},
                                {16'h1445, 16'h1449, 16'h144d, 16'h1451, 16'h1455, 16'h1459, 16'h145d, 16'h1461, 16'h1465, 16'h1469, 16'h146d, 16'h1471, 16'h1475, 16'h1479, 16'h147d, 16'h1481, 16'h1485, 16'h1489, 16'h148d, 16'h1491, 16'h1495, 16'h1499, 16'h149d, 16'h14a1, 16'h14a5, 16'h14a9, 16'h14ad, 16'h14b1, 16'h14b5, 16'h14b9, 16'h14bd, 16'h14c1, 16'h14c5, 16'h14c9, 16'h14cd, 16'h14d1, 16'h1553, 16'h155b, 16'h1563, 16'h156b, 16'h1573, 16'h157b, 16'h1583, 16'h158b, 16'h1593, 16'h159b, 16'h15a3, 16'h15ab, 16'h15b3, 16'h15bb, 16'h15c3, 16'h15cb, 16'h15d3, 16'h15db, 16'h15e3, 16'h15eb, 16'h15f3, 16'h15fb, 16'h1603, 16'h160b, 16'h1613, 16'h161b, 16'h1623, 16'h162b},
                                {16'h1633, 16'h163b, 16'h1643, 16'h164b, 16'h1653, 16'h165b, 16'h1663, 16'h166b, 16'h1673, 16'h167b, 16'h1683, 16'h168b, 16'h1693, 16'h169b, 16'h16a3, 16'h16ab, 16'h16b3, 16'h16bb, 16'h16c3, 16'h16cb, 16'h16d3, 16'h16db, 16'h16e3, 16'h16eb, 16'h16f3, 16'h16fb, 16'h1703, 16'h170b, 16'h1713, 16'h171b, 16'h1723, 16'h172b, 16'h1733, 16'h173b, 16'h1743, 16'h174b, 16'h1753, 16'h175b, 16'h1763, 16'h176b, 16'h1773, 16'h177b, 16'h1783, 16'h178b, 16'h1793, 16'h179b, 16'h17a3, 16'h17ab, 16'h17b3, 16'h17bb, 16'h17c3, 16'h17cb, 16'h17d3, 16'h17db, 16'h17e3, 16'h17eb, 16'h17f3, 16'h17fb, 16'h1803, 16'h180b, 16'h1813, 16'h181b, 16'h1823, 16'h182b},
                                {16'h1833, 16'h183b, 16'h1843, 16'h184b, 16'h1853, 16'h185b, 16'h1863, 16'h186b, 16'h1873, 16'h187b, 16'h1883, 16'h188b, 16'h1893, 16'h189b, 16'h18a3, 16'h18ab, 16'h18b3, 16'h18bb, 16'h18c3, 16'h18cb, 16'h18d3, 16'h18db, 16'h18e3, 16'h18eb, 16'h18f3, 16'h18fb, 16'h1903, 16'h190b, 16'h1913, 16'h191b, 16'h1923, 16'h192b, 16'h1933, 16'h193b, 16'h1943, 16'h194b, 16'h1953, 16'h195b, 16'h1963, 16'h196b, 16'h1973, 16'h197b, 16'h1983, 16'h198b, 16'h1993, 16'h199b, 16'h19a3, 16'h19ab, 16'h19b3, 16'h19bb, 16'h19c3, 16'h19cb, 16'h19d3, 16'h19db, 16'h19e3, 16'h19eb, 16'h19f3, 16'h19fb, 16'h1a03, 16'h1a0b, 16'h1a13, 16'h1a1b, 16'h1a23, 16'h1a2b},
                                {16'h1a33, 16'h1a3b, 16'h1a43, 16'h1a4b, 16'h1a53, 16'h1a5b, 16'h1a63, 16'h1a6b, 16'h1a73, 16'h1a7b, 16'h1a83, 16'h1a8b, 16'h1a93, 16'h1a9b, 16'h1aa3, 16'h1aab, 16'h1ab3, 16'h1abb, 16'h1ac3, 16'h1acb, 16'h1ad3, 16'h1adb, 16'h1ae3, 16'h1aeb, 16'h1af3, 16'h1afb, 16'h1b03, 16'h1b0b, 16'h1b13, 16'h1b1b, 16'h1b23, 16'h1b2b, 16'h1b33, 16'h1b3b, 16'h1b43, 16'h1b4b, 16'h1b53, 16'h1b5b, 16'h1b63, 16'h1b6b, 16'h1b73, 16'h1b7b, 16'h1b83, 16'h1b8b, 16'h1b93, 16'h1b9b, 16'h1ba3, 16'h1bab, 16'h1bb3, 16'h1bbb, 16'h1bc3, 16'h1bcb, 16'h1bd3, 16'h1bdb, 16'h1be3, 16'h1beb, 16'h1bf3, 16'h1bfb, 16'h1c03, 16'h1c0b, 16'h1c13, 16'h1c1b, 16'h1c23, 16'h1c2b},
                                {16'h1c33, 16'h1c3b, 16'h1c43, 16'h1c4b, 16'h1c53, 16'h1c5b, 16'h1c63, 16'h1c6b, 16'h1c73, 16'h1c7b, 16'h1c83, 16'h1c8b, 16'h1c93, 16'h1c9b, 16'h1ca3, 16'h1cab, 16'h1cb3, 16'h1cbb, 16'h1cc3, 16'h1ccb, 16'h1cd3, 16'h1cdb, 16'h1ce3, 16'h1ceb, 16'h1cf3, 16'h1cfb, 16'h1d03, 16'h1d0b, 16'h1d13, 16'h1d1b, 16'h1d23, 16'h1d2b, 16'h1d33, 16'h1d3b, 16'h1d43, 16'h1d4b, 16'h1d53, 16'h1d5b, 16'h1d63, 16'h1d6b, 16'h1d73, 16'h1d7b, 16'h1d83, 16'h1d8b, 16'h1d93, 16'h1d9b, 16'h1da3, 16'h1dab, 16'h1db3, 16'h1dbb, 16'h1dc3, 16'h1dcb, 16'h1dd3, 16'h1ddb, 16'h1de3, 16'h1deb, 16'h1df3, 16'h1dfb, 16'h1e03, 16'h1e0b, 16'h1e13, 16'h1e1b, 16'h1e23, 16'h1e2b},
                                {16'h1e33, 16'h1e3b, 16'h1e43, 16'h1e4b, 16'h1e53, 16'h1e5b, 16'h1e63, 16'h1e6b, 16'h1e73, 16'h1e7b, 16'h1e83, 16'h1e8b, 16'h1e93, 16'h1e9b, 16'h1ea3, 16'h1eab, 16'h1eb3, 16'h1ebb, 16'h1ec3, 16'h1ecb, 16'h1ed3, 16'h1edb, 16'h1ee3, 16'h1eeb, 16'h1ef3, 16'h1efb, 16'h1f03, 16'h1f0b, 16'h1f13, 16'h1f1b, 16'h1f23, 16'h1f2b, 16'h1f33, 16'h1f3b, 16'h1f43, 16'h1f4b, 16'h1f53, 16'h1f5b, 16'h1f63, 16'h1f6b, 16'h1f73, 16'h1f7b, 16'h1f83, 16'h1f8b, 16'h1f93, 16'h1f9b, 16'h1fa3, 16'h1fab, 16'h1fb3, 16'h1fbb, 16'h1fc3, 16'h1fcb, 16'h1fd3, 16'h1fdb, 16'h1fe3, 16'h1feb, 16'h1ff3, 16'h1ffb, 16'h2003, 16'h200b, 16'h2013, 16'h201b, 16'h2023, 16'h202b},
                                {16'h2033, 16'h203b, 16'h2043, 16'h204b, 16'h2053, 16'h205b, 16'h2063, 16'h206b, 16'h2073, 16'h207b, 16'h2083, 16'h208b, 16'h2093, 16'h209b, 16'h20a3, 16'h20ab, 16'h20b3, 16'h20bb, 16'h20c3, 16'h20cb, 16'h20d3, 16'h20db, 16'h20e3, 16'h20eb, 16'h20f3, 16'h20fb, 16'h2103, 16'h210b, 16'h2113, 16'h211b, 16'h2123, 16'h212b, 16'h2133, 16'h213b, 16'h2143, 16'h214b, 16'h2153, 16'h215b, 16'h2163, 16'h216b, 16'h2173, 16'h217b, 16'h2183, 16'h218b, 16'h2193, 16'h219b, 16'h21a3, 16'h21ab, 16'h21b3, 16'h21bb, 16'h21c3, 16'h21cb, 16'h21d3, 16'h21db, 16'h21e3, 16'h21eb, 16'h21f3, 16'h21fb, 16'h2203, 16'h220b, 16'h2213, 16'h221b, 16'h2223, 16'h222b},
                                {16'h2233, 16'h223b, 16'h2243, 16'h224b, 16'h2253, 16'h225b, 16'h2263, 16'h226b, 16'h2273, 16'h227b, 16'h2283, 16'h228b, 16'h2293, 16'h229b, 16'h22a3, 16'h22ab, 16'h22b3, 16'h22bb, 16'h22c3, 16'h22cb, 16'h22d3, 16'h22db, 16'h22e3, 16'h22eb, 16'h22f3, 16'h22fb, 16'h2303, 16'h230b, 16'h2313, 16'h231b, 16'h2323, 16'h232b, 16'h2333, 16'h233b, 16'h2343, 16'h234b, 16'h2353, 16'h235b, 16'h2363, 16'h236b, 16'h2373, 16'h237b, 16'h2383, 16'h238b, 16'h2393, 16'h239b, 16'h23a3, 16'h23ab, 16'h23b3, 16'h23bb, 16'h23c3, 16'h23cb, 16'h23d3, 16'h23db, 16'h23e3, 16'h23eb, 16'h23f3, 16'h23fb, 16'h2403, 16'h240b, 16'h2413, 16'h241b, 16'h2423, 16'h242b},
                                {16'h2433, 16'h243b, 16'h2443, 16'h244b, 16'h2453, 16'h245b, 16'h2463, 16'h246b, 16'h2473, 16'h247b, 16'h2483, 16'h248b, 16'h2493, 16'h249b, 16'h24a3, 16'h24ab, 16'h24b3, 16'h24bb, 16'h24c3, 16'h24cb, 16'h24d3, 16'h24db, 16'h24e3, 16'h24eb, 16'h24f3, 16'h24fb, 16'h2503, 16'h250b, 16'h2513, 16'h251b, 16'h2523, 16'h252b, 16'h2533, 16'h253b, 16'h2543, 16'h254b, 16'h2553, 16'h255b, 16'h2563, 16'h256b, 16'h2573, 16'h257b, 16'h2583, 16'h258b, 16'h2593, 16'h259b, 16'h25a3, 16'h25ab, 16'h25b3, 16'h25bb, 16'h25c3, 16'h25cb, 16'h25d3, 16'h25db, 16'h25e3, 16'h25eb, 16'h25f3, 16'h25fb, 16'h2603, 16'h260b, 16'h2613, 16'h261b, 16'h2623, 16'h262b},
                                {16'h2633, 16'h263b, 16'h2643, 16'h264b, 16'h2653, 16'h265b, 16'h2663, 16'h266b, 16'h2673, 16'h267b, 16'h2683, 16'h268b, 16'h2693, 16'h269b, 16'h26a3, 16'h26ab, 16'h26b3, 16'h26bb, 16'h26c3, 16'h26cb, 16'h26d3, 16'h26db, 16'h26e3, 16'h26eb, 16'h26f3, 16'h26fb, 16'h2703, 16'h270b, 16'h2713, 16'h271b, 16'h2723, 16'h272b, 16'h2733, 16'h273b, 16'h2743, 16'h274b, 16'h2753, 16'h275b, 16'h2763, 16'h276b, 16'h2773, 16'h277b, 16'h2783, 16'h278b, 16'h2793, 16'h279b, 16'h27a3, 16'h27ab, 16'h27b3, 16'h27bb, 16'h27c3, 16'h27cb, 16'h27d3, 16'h27db, 16'h27e3, 16'h27eb, 16'h27f3, 16'h27fb, 16'h2803, 16'h280b, 16'h2813, 16'h281b, 16'h2823, 16'h282b},
                                {16'h2833, 16'h283b, 16'h2843, 16'h284b, 16'h2853, 16'h285b, 16'h2863, 16'h286b, 16'h2873, 16'h287b, 16'h2883, 16'h288b, 16'h2893, 16'h289b, 16'h28a3, 16'h28ab, 16'h28b3, 16'h28bb, 16'h28c3, 16'h28cb, 16'h28d3, 16'h28db, 16'h28e3, 16'h28eb, 16'h28f3, 16'h28fb, 16'h2903, 16'h290b, 16'h2913, 16'h291b, 16'h2923, 16'h292b, 16'h2933, 16'h293b, 16'h2943, 16'h294b, 16'h2953, 16'h295b, 16'h2963, 16'h296b, 16'h2973, 16'h297b, 16'h2983, 16'h298b, 16'h2993, 16'h299b, 16'h29a3, 16'h29ab, 16'h29b3, 16'h29bb, 16'h29c3, 16'h29cb, 16'h29d3, 16'h29db, 16'h29e3, 16'h29eb, 16'h29f3, 16'h29fb, 16'h2a03, 16'h2a0b, 16'h2a13, 16'h2a1b, 16'h2a23, 16'h2a2b},
                                {16'h2a33, 16'h2a3b, 16'h2a43, 16'h2a4b, 16'h2a53, 16'h2a5b, 16'h2a63, 16'h2a6b, 16'h2a73, 16'h2a7b, 16'h2a83, 16'h2a8b, 16'h2a93, 16'h2a9b, 16'h2aa3, 16'h2aab, 16'h2ab3, 16'h2abb, 16'h2ac3, 16'h2acb, 16'h2ad3, 16'h2adb, 16'h2ae3, 16'h2aeb, 16'h2af3, 16'h2afb, 16'h2b03, 16'h2b0b, 16'h2b13, 16'h2b1b, 16'h2b23, 16'h2b2b, 16'h2b33, 16'h2b3b, 16'h2b43, 16'h2b4b, 16'h2b53, 16'h2b5b, 16'h2b63, 16'h2b6b, 16'h2b73, 16'h2b7b, 16'h2b83, 16'h2b8b, 16'h2b93, 16'h2b9b, 16'h2ba3, 16'h2ba3, 16'h2ba3, 16'h2ba3, 16'h2ba3, 16'h2ba3, 16'h2ba3, 16'h2ba3, 16'h2ba3, 16'h2ba3, 16'h2ba3, 16'h2ba3, 16'h2ba3, 16'h2baa, 16'h2bb2, 16'h2bba, 16'h2bc2, 16'h2bca},
                                {16'h2bd2, 16'h2bda, 16'h2be2, 16'h2bea, 16'h2bf2, 16'h2bfa, 16'h2c02, 16'h2c0a, 16'h2c12, 16'h2c1a, 16'h2c22, 16'h2c2a, 16'h2c32, 16'h2c3a, 16'h2c42, 16'h2c4a, 16'h2c52, 16'h2c5a, 16'h2c62, 16'h2c6a, 16'h2c72, 16'h2c7a, 16'h2c82, 16'h2c8a, 16'h2c92, 16'h2c9a, 16'h2ca2, 16'h2caa, 16'h2cb2, 16'h2cba, 16'h2cc2, 16'h2cca, 16'h2cd2, 16'h2cda, 16'h2ce2, 16'h2cea, 16'h2cf2, 16'h2cfa, 16'h2d02, 16'h2d0a, 16'h2d12, 16'h2d1a, 16'h2d22, 16'h2d2a, 16'h2d32, 16'h2d3a, 16'h2d42, 16'h2d4a, 16'h2d52, 16'h2d5a, 16'h2d62, 16'h2d6a, 16'h2d72, 16'h2d7a, 16'h2d82, 16'h2d8a, 16'h2d92, 16'h2d9a, 16'h2da2, 16'h2daa, 16'h2db2, 16'h2dba, 16'h2dc2, 16'h2dca},
                                {16'h2dd2, 16'h2dda, 16'h2de2, 16'h2dea, 16'h2df2, 16'h2dfa, 16'h2e02, 16'h2e0a, 16'h2e12, 16'h2e1a, 16'h2e22, 16'h2e2a, 16'h2e32, 16'h2e3a, 16'h2e42, 16'h2e4a, 16'h2e52, 16'h2e5a, 16'h2e62, 16'h2e6a, 16'h2e72, 16'h2e7a, 16'h2e82, 16'h2e8a, 16'h2e92, 16'h2e9a, 16'h2ea2, 16'h2eaa, 16'h2eb2, 16'h2eba, 16'h2ec2, 16'h2eca, 16'h2ed2, 16'h2eda, 16'h2ee2, 16'h2eea, 16'h2ef2, 16'h2efa, 16'h2f02, 16'h2f0a, 16'h2f12, 16'h2f1a, 16'h2f22, 16'h2f2a, 16'h2f32, 16'h2f3a, 16'h2f42, 16'h2f4a, 16'h2f52, 16'h2f5a, 16'h2f62, 16'h2f6a, 16'h2f72, 16'h2f7a, 16'h2f82, 16'h2f8a, 16'h2f92, 16'h2f9a, 16'h2fa2, 16'h2faa, 16'h2fb2, 16'h2fba, 16'h2fc2, 16'h2fca},
                                {16'h2fd2, 16'h2fda, 16'h2fe2, 16'h2fea, 16'h2ff2, 16'h2ffa, 16'h3002, 16'h300a, 16'h3012, 16'h301a, 16'h3022, 16'h302a, 16'h3032, 16'h303a, 16'h3042, 16'h304a, 16'h3052, 16'h305a, 16'h3062, 16'h306a, 16'h3072, 16'h307a, 16'h3082, 16'h308a, 16'h3092, 16'h309a, 16'h30a2, 16'h30aa, 16'h30b2, 16'h30ba, 16'h30c2, 16'h30ca, 16'h30d2, 16'h30da, 16'h30e2, 16'h30ea, 16'h30f2, 16'h30fa, 16'h3102, 16'h310a, 16'h3112, 16'h311a, 16'h3122, 16'h312a, 16'h3132, 16'h313a, 16'h3142, 16'h314a, 16'h3152, 16'h315a, 16'h3162, 16'h316a, 16'h3172, 16'h317a, 16'h3182, 16'h318a, 16'h3192, 16'h319a, 16'h31a2, 16'h31aa, 16'h31b2, 16'h31ba, 16'h31c2, 16'h31ca},
                                {16'h31d2, 16'h31da, 16'h31e2, 16'h31ea, 16'h31f2, 16'h31fa, 16'h3202, 16'h320a, 16'h3212, 16'h321a, 16'h3222, 16'h322a, 16'h3232, 16'h323a, 16'h3242, 16'h324a, 16'h3252, 16'h325a, 16'h3262, 16'h326a, 16'h3272, 16'h327a, 16'h3282, 16'h328a, 16'h3292, 16'h329a, 16'h32a2, 16'h32aa, 16'h32b2, 16'h32ba, 16'h32c2, 16'h32ca, 16'h32d2, 16'h32da, 16'h32e2, 16'h32ea, 16'h32f2, 16'h32fa, 16'h3302, 16'h330a, 16'h3312, 16'h331a, 16'h3322, 16'h332a, 16'h3332, 16'h333a, 16'h3342, 16'h334a, 16'h3352, 16'h335a, 16'h3362, 16'h336a, 16'h3372, 16'h337a, 16'h3382, 16'h338a, 16'h3392, 16'h339a, 16'h33a2, 16'h33aa, 16'h33b2, 16'h33ba, 16'h33c2, 16'h33ca},
                                {16'h33d2, 16'h33da, 16'h33e2, 16'h33ea, 16'h33f2, 16'h33fa, 16'h3402, 16'h340a, 16'h3412, 16'h341a, 16'h3422, 16'h342a, 16'h3432, 16'h343a, 16'h3442, 16'h344a, 16'h3452, 16'h345a, 16'h3462, 16'h346a, 16'h3472, 16'h347a, 16'h3482, 16'h348a, 16'h3492, 16'h349a, 16'h34a2, 16'h34aa, 16'h34b2, 16'h34ba, 16'h34c2, 16'h34ca, 16'h34d2, 16'h34da, 16'h34e2, 16'h34ea, 16'h34f2, 16'h34fa, 16'h3502, 16'h350a, 16'h3512, 16'h351a, 16'h3522, 16'h352a, 16'h3532, 16'h353a, 16'h3542, 16'h354a, 16'h3552, 16'h355a, 16'h3562, 16'h356a, 16'h3572, 16'h357a, 16'h3582, 16'h358a, 16'h3592, 16'h359a, 16'h35a2, 16'h35aa, 16'h35b2, 16'h35ba, 16'h35c2, 16'h35ca},
                                {16'h35d2, 16'h35da, 16'h360f, 16'h3617, 16'h361f, 16'h3627, 16'h362f, 16'h3637, 16'h363f, 16'h3647, 16'h364f, 16'h3657, 16'h365f, 16'h3667, 16'h366f, 16'h3677, 16'h367f, 16'h3687, 16'h368f, 16'h3697, 16'h369f, 16'h36a7, 16'h36af, 16'h36b7, 16'h36bf, 16'h36c7, 16'h36cf, 16'h36d7, 16'h36df, 16'h36e7, 16'h36ef, 16'h36f7, 16'h36ff, 16'h3707, 16'h370f, 16'h3717, 16'h371f, 16'h3727, 16'h372f, 16'h3737, 16'h373f, 16'h3747, 16'h374f, 16'h3757, 16'h375f, 16'h3767, 16'h376f, 16'h3777, 16'h377f, 16'h3787, 16'h378f, 16'h3797, 16'h379f, 16'h37a7, 16'h37af, 16'h37b7, 16'h37bf, 16'h37c7, 16'h37cf, 16'h37d7, 16'h37df, 16'h37e7, 16'h37ef, 16'h37f7},
                                {16'h37ff, 16'h3807, 16'h380f, 16'h3817, 16'h381f, 16'h3827, 16'h382f, 16'h3837, 16'h383f, 16'h3847, 16'h384f, 16'h3857, 16'h385f, 16'h3867, 16'h386f, 16'h3877, 16'h387f, 16'h3887, 16'h388f, 16'h3897, 16'h389f, 16'h38a7, 16'h38af, 16'h38b7, 16'h38bf, 16'h38c7, 16'h38cf, 16'h38d7, 16'h38df, 16'h38e7, 16'h38ef, 16'h38f7, 16'h38ff, 16'h3907, 16'h390f, 16'h3917, 16'h391f, 16'h3927, 16'h392f, 16'h3937, 16'h393f, 16'h3947, 16'h394f, 16'h3957, 16'h395f, 16'h3967, 16'h396f, 16'h3977, 16'h397f, 16'h3987, 16'h398f, 16'h3997, 16'h399f, 16'h39a7, 16'h39af, 16'h39b7, 16'h39bf, 16'h39c7, 16'h39cf, 16'h39d7, 16'h39df, 16'h39e7, 16'h39ef, 16'h39f7},
                                {16'h39ff, 16'h3a07, 16'h3a0f, 16'h3a17, 16'h3a1f, 16'h3a27, 16'h3a2f, 16'h3a37, 16'h3a3f, 16'h3a47, 16'h3a4f, 16'h3a57, 16'h3a5f, 16'h3a67, 16'h3a6f, 16'h3a77, 16'h3a7f, 16'h3a87, 16'h3a8f, 16'h3a97, 16'h3a9f, 16'h3aa7, 16'h3aaf, 16'h3ab7, 16'h3abf, 16'h3ac7, 16'h3acf, 16'h3ad7, 16'h3adf, 16'h3ae7, 16'h3aef, 16'h3af7, 16'h3aff, 16'h3b07, 16'h3b0f, 16'h3b17, 16'h3b1f, 16'h3b27, 16'h3b2f, 16'h3b37, 16'h3b3f, 16'h3b47, 16'h3b4f, 16'h3b57, 16'h3b5f, 16'h3b67, 16'h3b6f, 16'h3b77, 16'h3b7f, 16'h3b87, 16'h3b8f, 16'h3b97, 16'h3b9f, 16'h3ba7, 16'h3baf, 16'h3bb7, 16'h3bbf, 16'h3bc7, 16'h3bcf, 16'h3bd7, 16'h3bdf, 16'h3be7, 16'h3bef, 16'h3bf7},
                                {16'h3bff, 16'h3c07, 16'h3c0f, 16'h3c17, 16'h3c1f, 16'h3c27, 16'h3c2f, 16'h3c37, 16'h3c3f, 16'h3c47, 16'h3c4f, 16'h3c57, 16'h3c5f, 16'h3c67, 16'h3c6f, 16'h3c77, 16'h3c7f, 16'h3c87, 16'h3c8f, 16'h3c97, 16'h3c9f, 16'h3ca7, 16'h3caf, 16'h3cb7, 16'h3cbf, 16'h3cc7, 16'h3ccf, 16'h3cd7, 16'h3cdf, 16'h3ce7, 16'h3cef, 16'h3cf7, 16'h3cff, 16'h3d07, 16'h3d0f, 16'h3d17, 16'h3d1f, 16'h3d27, 16'h3d2f, 16'h3d37, 16'h3d3f, 16'h3d47, 16'h3d4f, 16'h3d57, 16'h3d5f, 16'h3d67, 16'h3d6f, 16'h3d77, 16'h3d7f, 16'h3d87, 16'h3d8f, 16'h3d97, 16'h3d9f, 16'h3da7, 16'h3daf, 16'h3db7, 16'h3dbf, 16'h3dc7, 16'h3dcf, 16'h3dd7, 16'h3ddf, 16'h3de7, 16'h3def, 16'h3df7},
                                {16'h3dff, 16'h3e07, 16'h3e0f, 16'h3e17, 16'h3e1f, 16'h3e27, 16'h3e2f, 16'h3e37, 16'h3e3f, 16'h3e47, 16'h3e4f, 16'h3e57, 16'h3e5f, 16'h3e67, 16'h3e6f, 16'h3e77, 16'h3e7f, 16'h3e87, 16'h3e8f, 16'h3e97, 16'h3e9f, 16'h3ea7, 16'h3eaf, 16'h3eb7, 16'h3ebf, 16'h3ec7, 16'h3ecf, 16'h3ed7, 16'h3edf, 16'h3ee7, 16'h3eef, 16'h3ef7, 16'h3eff, 16'h3f07, 16'h3f0f, 16'h3f17, 16'h3f1f, 16'h3f27, 16'h3f2f, 16'h3f37, 16'h3f3f, 16'h3f47, 16'h3f4f, 16'h3f57, 16'h3f5f, 16'h3f67, 16'h3f6f, 16'h3f77, 16'h3f7f, 16'h3f87, 16'h3f8f, 16'h3f97, 16'h3f9f, 16'h3fa7, 16'h3faf, 16'h3fb7, 16'h3fbf, 16'h3fc7, 16'h3fcf, 16'h3fd7, 16'h3fdf, 16'h3fe7, 16'h3fef, 16'h3ff7},
                                {16'h3fff, 16'h3fbb, 16'h3fab, 16'h3f9b, 16'h3f8b, 16'h3f7b, 16'h3f6b, 16'h3f5b, 16'h3f4b, 16'h3f3b, 16'h3f2b, 16'h3f1b, 16'h3f0b, 16'h3efb, 16'h3eeb, 16'h3edb, 16'h3ecb, 16'h3ebb, 16'h3eab, 16'h3e9b, 16'h3e8b, 16'h3e7b, 16'h3e6b, 16'h3e5b, 16'h3e4b, 16'h3e3b, 16'h3e2b, 16'h3e1b, 16'h3e0b, 16'h3dfb, 16'h3deb, 16'h3ddb, 16'h3dcb, 16'h3dbb, 16'h3dab, 16'h3d9b, 16'h3d8b, 16'h3d7b, 16'h3d6b, 16'h3d5b, 16'h3d4b, 16'h3d3b, 16'h3d2b, 16'h3d1b, 16'h3d0b, 16'h3cfb, 16'h3ceb, 16'h3cdb, 16'h3ccb, 16'h3cbb, 16'h3cab, 16'h3c9b, 16'h3c8b, 16'h3c7b, 16'h3c6b, 16'h3c5b, 16'h3c4b, 16'h3c3b, 16'h3c2b, 16'h3c1b, 16'h3c0b, 16'h3bfb, 16'h3beb, 16'h3bdb},
                                {16'h3bcb, 16'h3bbb, 16'h3bab, 16'h3b9b, 16'h3b8b, 16'h3b7b, 16'h3b6b, 16'h3b5b, 16'h3b4b, 16'h3b3b, 16'h3b2b, 16'h3b1b, 16'h3b0b, 16'h3afb, 16'h3aeb, 16'h3adb, 16'h3acb, 16'h3abb, 16'h3aab, 16'h3a9b, 16'h3a8b, 16'h3a7b, 16'h3a6b, 16'h3a5b, 16'h3a4b, 16'h3a3b, 16'h3a2b, 16'h3a1b, 16'h3a0b, 16'h39fb, 16'h39eb, 16'h39db, 16'h39cb, 16'h39bb, 16'h39ab, 16'h399b, 16'h398b, 16'h397b, 16'h396b, 16'h395b, 16'h394b, 16'h393b, 16'h392b, 16'h391b, 16'h390b, 16'h38fb, 16'h38eb, 16'h38db, 16'h38cb, 16'h38bb, 16'h38ab, 16'h389b, 16'h388b, 16'h387b, 16'h386b, 16'h385b, 16'h384b, 16'h383b, 16'h382b, 16'h381b, 16'h380b, 16'h37fb, 16'h37eb, 16'h37db},
                                {16'h37cb, 16'h37bb, 16'h37ab, 16'h379b, 16'h378b, 16'h377b, 16'h376b, 16'h375b, 16'h374b, 16'h373b, 16'h372b, 16'h371b, 16'h370b, 16'h36fb, 16'h36eb, 16'h36db, 16'h36cb, 16'h36bb, 16'h36ab, 16'h369b, 16'h368b, 16'h367b, 16'h366b, 16'h365b, 16'h364b, 16'h363b, 16'h362b, 16'h361b, 16'h360b, 16'h35fb, 16'h35eb, 16'h35db, 16'h35cb, 16'h35bb, 16'h35ab, 16'h359b, 16'h358b, 16'h357b, 16'h356b, 16'h355b, 16'h354b, 16'h353b, 16'h352b, 16'h351b, 16'h350b, 16'h34fb, 16'h34eb, 16'h34db, 16'h34cb, 16'h34bb, 16'h34ab, 16'h349b, 16'h348b, 16'h347b, 16'h346b, 16'h345b, 16'h344b, 16'h343b, 16'h342b, 16'h341b, 16'h340b, 16'h33fb, 16'h33eb, 16'h33db},
                                {16'h33cb, 16'h33bb, 16'h33ab, 16'h339b, 16'h338b, 16'h337b, 16'h336b, 16'h335b, 16'h334b, 16'h333b, 16'h332b, 16'h331b, 16'h330b, 16'h32fb, 16'h32eb, 16'h32db, 16'h32db, 16'h32db, 16'h32db, 16'h32db, 16'h32db, 16'h32db, 16'h32db, 16'h32db, 16'h32db, 16'h32db, 16'h32db, 16'h32db, 16'h32db, 16'h32db, 16'h32db, 16'h32db, 16'h32db, 16'h32db, 16'h32db, 16'h32db, 16'h32db, 16'h32db, 16'h32db, 16'h32db, 16'h32db, 16'h32db, 16'h32db, 16'h32db, 16'h32d9, 16'h32d6, 16'h32d3, 16'h32d0, 16'h32cd, 16'h32ca, 16'h32c7, 16'h32c4, 16'h32c1, 16'h32be, 16'h32bb, 16'h32b8, 16'h32b5, 16'h32b2, 16'h32af, 16'h32ac, 16'h32a9, 16'h32a6, 16'h32a3, 16'h32a0},
                                {16'h329d, 16'h329a, 16'h3297, 16'h3294, 16'h3291, 16'h328e, 16'h328b, 16'h3288, 16'h3285, 16'h3282, 16'h327f, 16'h327c, 16'h3279, 16'h3276, 16'h3273, 16'h3270, 16'h326d, 16'h326a, 16'h3267, 16'h3264, 16'h3261, 16'h325e, 16'h325b, 16'h3258, 16'h3255, 16'h3252, 16'h324f, 16'h324c, 16'h3249, 16'h3246, 16'h3243, 16'h3240, 16'h323d, 16'h323a, 16'h3237, 16'h3234, 16'h3231, 16'h322e, 16'h322b, 16'h3228, 16'h3225, 16'h3222, 16'h321f, 16'h321c, 16'h3219, 16'h3216, 16'h3213, 16'h3210, 16'h320d, 16'h320a, 16'h3207, 16'h3204, 16'h3201, 16'h31fe, 16'h31fb, 16'h31f8, 16'h31f5, 16'h31f2, 16'h31ef, 16'h31ec, 16'h31e9, 16'h31e6, 16'h31e3, 16'h31e0},
                                {16'h31dd, 16'h31da, 16'h31d7, 16'h31d4, 16'h31d1, 16'h31ce, 16'h31cb, 16'h31c8, 16'h31c5, 16'h31c2, 16'h31bf, 16'h31bc, 16'h31b9, 16'h31b6, 16'h31b3, 16'h31b0, 16'h31ad, 16'h31aa, 16'h31a7, 16'h31a4, 16'h31a1, 16'h319e, 16'h319b, 16'h3198, 16'h3195, 16'h3192, 16'h318f, 16'h318c, 16'h3189, 16'h3186, 16'h3183, 16'h3180, 16'h317d, 16'h317a, 16'h3177, 16'h3174, 16'h3171, 16'h316e, 16'h316b, 16'h3168, 16'h3165, 16'h3162, 16'h315f, 16'h315c, 16'h3159, 16'h3156, 16'h3153, 16'h3150, 16'h314d, 16'h314a, 16'h3147, 16'h3144, 16'h3141, 16'h313e, 16'h313b, 16'h3138, 16'h3135, 16'h3132, 16'h312f, 16'h312c, 16'h3129, 16'h3126, 16'h3123, 16'h3120},
                                {16'h311d, 16'h311a, 16'h3117, 16'h3114, 16'h3111, 16'h310e, 16'h310b, 16'h3108, 16'h3105, 16'h3102, 16'h30ff, 16'h30fc, 16'h30f9, 16'h30f6, 16'h30f3, 16'h30f0, 16'h30ed, 16'h30ea, 16'h30e7, 16'h30e4, 16'h30e1, 16'h30de, 16'h30db, 16'h30d8, 16'h30d5, 16'h30d2, 16'h30cf, 16'h30cc, 16'h30c9, 16'h30c6, 16'h30c3, 16'h30c0, 16'h30bd, 16'h30ba, 16'h30b7, 16'h30b4, 16'h30b1, 16'h30ae, 16'h30ab, 16'h30a8, 16'h30a5, 16'h30a2, 16'h309f, 16'h309c, 16'h3099, 16'h3096, 16'h3093, 16'h3090, 16'h308d, 16'h308a, 16'h3087, 16'h3084, 16'h3081, 16'h307e, 16'h307b, 16'h3078, 16'h3075, 16'h3072, 16'h306f, 16'h306c, 16'h3069, 16'h3066, 16'h3063, 16'h3060},
                                {16'h305d, 16'h305a, 16'h3057, 16'h3054, 16'h3051, 16'h304e, 16'h304b, 16'h3048, 16'h3045, 16'h3042, 16'h303f, 16'h303c, 16'h3039, 16'h3036, 16'h3033, 16'h3030, 16'h302d, 16'h302a, 16'h3027, 16'h3024, 16'h3021, 16'h301e, 16'h301b, 16'h3018, 16'h3015, 16'h3012, 16'h300f, 16'h300c, 16'h3009, 16'h3006, 16'h3003, 16'h3000, 16'h2ffd, 16'h2ffa, 16'h2ff7, 16'h2ff4, 16'h2ff1, 16'h2fee, 16'h2feb, 16'h2fe8, 16'h2fe5, 16'h2fe2, 16'h2fdf, 16'h2fdc, 16'h2fd9, 16'h2fd6, 16'h2fd3, 16'h2fd0, 16'h2fcd, 16'h2fca, 16'h2fc7, 16'h2fc4, 16'h2fc1, 16'h2fbe, 16'h2fbb, 16'h2fb8, 16'h2fb5, 16'h2fb2, 16'h2faf, 16'h2fac, 16'h2fa9, 16'h2fa6, 16'h2fa3, 16'h2fa0},
                                {16'h2f9d, 16'h2f9a, 16'h2f97, 16'h2f94, 16'h2f91, 16'h2f8e, 16'h2f8b, 16'h2f88, 16'h2f85, 16'h2f82, 16'h2f7f, 16'h2f7c, 16'h2f79, 16'h2f76, 16'h2f73, 16'h2f70, 16'h2f6d, 16'h2f6a, 16'h2f67, 16'h2f64, 16'h2f61, 16'h2f5e, 16'h2f5b, 16'h2f58, 16'h2f55, 16'h2f52, 16'h2f4f, 16'h2f4c, 16'h2f49, 16'h2f46, 16'h2f43, 16'h2f40, 16'h2f3d, 16'h2f3a, 16'h2f37, 16'h2f34, 16'h2f31, 16'h2f2e, 16'h2f2b, 16'h2f28, 16'h2f25, 16'h2f22, 16'h2f1f, 16'h2f1c, 16'h2f19, 16'h2f16, 16'h2f13, 16'h2f10, 16'h2f0d, 16'h2f0a, 16'h2f07, 16'h2f04, 16'h2f01, 16'h2efe, 16'h2efb, 16'h2ef8, 16'h2ef5, 16'h2ef2, 16'h2eef, 16'h2eec, 16'h2ee9, 16'h2ee6, 16'h2ee3, 16'h2ee0},
                                {16'h2edd, 16'h2eda, 16'h2ed7, 16'h2ed4, 16'h2ed1, 16'h2ece, 16'h2ecb, 16'h2ec8, 16'h2ec5, 16'h2ec2, 16'h2ebf, 16'h2ebc, 16'h2eb9, 16'h2eb6, 16'h2eb3, 16'h2eb0, 16'h2ead, 16'h2eaa, 16'h2ea7, 16'h2ea4, 16'h2ea1, 16'h2e9e, 16'h2e9b, 16'h2e98, 16'h2e95, 16'h2e92, 16'h2e8f, 16'h2e8c, 16'h2e89, 16'h2e86, 16'h2e83, 16'h2e80, 16'h2e7d, 16'h2e7a, 16'h2e77, 16'h2e74, 16'h2e71, 16'h2e6e, 16'h2e6b, 16'h2e68, 16'h2e65, 16'h2e62, 16'h2e5f, 16'h2e5c, 16'h2e59, 16'h2e56, 16'h2e53, 16'h2e50, 16'h2e4d, 16'h2e4a, 16'h2e47, 16'h2e44, 16'h2e41, 16'h2e3e, 16'h2e3b, 16'h2e38, 16'h2e35, 16'h2e32, 16'h2e2f, 16'h2e2c, 16'h2e29, 16'h2e26, 16'h2e23, 16'h2e20},
                                {16'h2e1d, 16'h2e1a, 16'h2e17, 16'h2e14, 16'h2e11, 16'h2e0e, 16'h2e0b, 16'h2e08, 16'h2e05, 16'h2e02, 16'h2dff, 16'h2dfc, 16'h2df9, 16'h2df6, 16'h2df3, 16'h2df0, 16'h2ded, 16'h2dea, 16'h2de7, 16'h2de4, 16'h2de1, 16'h2dde, 16'h2ddb, 16'h2dd8, 16'h2dd5, 16'h2dd2, 16'h2dcf, 16'h2dcc, 16'h2dc9, 16'h2dc6, 16'h2dc3, 16'h2dc0, 16'h2dbd, 16'h2dba, 16'h2db7, 16'h2db4, 16'h2db1, 16'h2dae, 16'h2dab, 16'h2da8, 16'h2da5, 16'h2da2, 16'h2d9f, 16'h2d9c, 16'h2d99, 16'h2d96, 16'h2d93, 16'h2d90, 16'h2d8d, 16'h2d8a, 16'h2d87, 16'h2d84, 16'h2d81, 16'h2d7e, 16'h2d7b, 16'h2d78, 16'h2d75, 16'h2d72, 16'h2d6f, 16'h2d6c, 16'h2d69, 16'h2d66, 16'h2d63, 16'h2d60},
                                {16'h2d5d, 16'h2d5a, 16'h2d57, 16'h2d54, 16'h2d51, 16'h2d4e, 16'h2d4b, 16'h2d48, 16'h2d45, 16'h2d42, 16'h2d3f, 16'h2d3c, 16'h2d39, 16'h2d36, 16'h2d33, 16'h2d30, 16'h2d2d, 16'h2d2a, 16'h2d27, 16'h2d24, 16'h2d21, 16'h2d1e, 16'h2d1b, 16'h2d18, 16'h2d15, 16'h2d12, 16'h2d0f, 16'h2d0c, 16'h2d09, 16'h2d06, 16'h2d03, 16'h2d00, 16'h2cfd, 16'h2cfa, 16'h2cf7, 16'h2cf4, 16'h2cf1, 16'h2cee, 16'h2ceb, 16'h2ce8, 16'h2ce5, 16'h2ce2, 16'h2cdf, 16'h2cdc, 16'h2cd9, 16'h2cd6, 16'h2cd3, 16'h2cd0, 16'h2ccd, 16'h2cca, 16'h2cca, 16'h2cca, 16'h2cca, 16'h2cca, 16'h2cca, 16'h2cca, 16'h2cca, 16'h2cca, 16'h2cca, 16'h2cca, 16'h2cca, 16'h2cca, 16'h2cca, 16'h2cca},
                                {16'h2cca, 16'h2cc9, 16'h2cc6, 16'h2cc3, 16'h2cc0, 16'h2cbd, 16'h2cba, 16'h2cb7, 16'h2cb4, 16'h2cb1, 16'h2cae, 16'h2cab, 16'h2ca8, 16'h2ca5, 16'h2ca2, 16'h2c9f, 16'h2c9c, 16'h2c99, 16'h2c96, 16'h2c93, 16'h2c90, 16'h2c8d, 16'h2c8a, 16'h2c87, 16'h2c84, 16'h2c81, 16'h2c7e, 16'h2c7b, 16'h2c78, 16'h2c75, 16'h2c72, 16'h2c6f, 16'h2c6c, 16'h2c69, 16'h2c66, 16'h2c63, 16'h2c60, 16'h2c5d, 16'h2c5a, 16'h2c57, 16'h2c54, 16'h2c51, 16'h2c4e, 16'h2c4b, 16'h2c48, 16'h2c45, 16'h2c42, 16'h2c3f, 16'h2c3c, 16'h2c39, 16'h2c36, 16'h2c33, 16'h2c30, 16'h2c2d, 16'h2c2a, 16'h2c27, 16'h2c24, 16'h2c21, 16'h2c1e, 16'h2c1b, 16'h2c18, 16'h2c15, 16'h2c12, 16'h2c0f},
                                {16'h2c0c, 16'h2c09, 16'h2c06, 16'h2c03, 16'h2c00, 16'h2bfd, 16'h2bfa, 16'h2bf7, 16'h2bf4, 16'h2bf1, 16'h2bee, 16'h2beb, 16'h2be8, 16'h2be5, 16'h2be2, 16'h2bdf, 16'h2bdc, 16'h2bd9, 16'h2bd6, 16'h2bd3, 16'h2bd0, 16'h2bcd, 16'h2bca, 16'h2bc7, 16'h2bc4, 16'h2bc1, 16'h2bbe, 16'h2bbb, 16'h2bb8, 16'h2bb5, 16'h2bb2, 16'h2baf, 16'h2bac, 16'h2ba9, 16'h2ba6, 16'h2ba3, 16'h2ba0, 16'h2b9d, 16'h2b9a, 16'h2b97, 16'h2b94, 16'h2b91, 16'h2b8e, 16'h2b8b, 16'h2b88, 16'h2b85, 16'h2b82, 16'h2b7f, 16'h2b7c, 16'h2b79, 16'h2b76, 16'h2b73, 16'h2b70, 16'h2b6d, 16'h2b6a, 16'h2b67, 16'h2b64, 16'h2b61, 16'h2b5e, 16'h2b5b, 16'h2b58, 16'h2b55, 16'h2b52, 16'h2b4f},
                                {16'h2b4c, 16'h2b49, 16'h2b46, 16'h2b43, 16'h2b40, 16'h2b3d, 16'h2b3a, 16'h2b37, 16'h2b34, 16'h2b31, 16'h2b2e, 16'h2b2b, 16'h2b28, 16'h2b25, 16'h2b22, 16'h2b1f, 16'h2b1c, 16'h2b19, 16'h2b16, 16'h2b13, 16'h2b10, 16'h2b0d, 16'h2b0a, 16'h2b07, 16'h2b04, 16'h2b01, 16'h2afe, 16'h2afb, 16'h2af8, 16'h2af5, 16'h2af2, 16'h2aef, 16'h2aec, 16'h2ae9, 16'h2ae6, 16'h2ae3, 16'h2ae0, 16'h2add, 16'h2ada, 16'h2ad7, 16'h2ad4, 16'h2ad1, 16'h2ace, 16'h2acb, 16'h2ac8, 16'h2ac5, 16'h2ac2, 16'h2abf, 16'h2abc, 16'h2ab9, 16'h2ab6, 16'h2ab3, 16'h2ab0, 16'h2aad, 16'h2aaa, 16'h2aa7, 16'h2aa4, 16'h2aa1, 16'h2a9e, 16'h2a9b, 16'h2a98, 16'h2a95, 16'h2a92, 16'h2a8f},
                                {16'h2a8c, 16'h2a89, 16'h2a86, 16'h2a83, 16'h2a80, 16'h2a7d, 16'h2a7a, 16'h2a77, 16'h2a74, 16'h2a71, 16'h2a6e, 16'h2a6b, 16'h2a68, 16'h2a65, 16'h2a62, 16'h2a5f, 16'h2a5c, 16'h2a59, 16'h2a56, 16'h2a53, 16'h2a50, 16'h2a4d, 16'h2a4a, 16'h2a47, 16'h2a44, 16'h2a41, 16'h2a3e, 16'h2a3b, 16'h2a38, 16'h2a35, 16'h2a32, 16'h2a2f, 16'h2a2c, 16'h2a29, 16'h2a26, 16'h2a23, 16'h2a20, 16'h2a1d, 16'h2a1a, 16'h2a17, 16'h2a14, 16'h2a11, 16'h2a0e, 16'h2a0b, 16'h2a08, 16'h2a05, 16'h2a02, 16'h29ff, 16'h29fc, 16'h29f9, 16'h29f6, 16'h29f3, 16'h29f0, 16'h29ed, 16'h29ea, 16'h29e7, 16'h29e4, 16'h29e1, 16'h29de, 16'h29db, 16'h29d8, 16'h29d5, 16'h29d2, 16'h29cf},
                                {16'h29cc, 16'h29c9, 16'h29c6, 16'h29c3, 16'h29c0, 16'h29bd, 16'h29ba, 16'h29b7, 16'h29b4, 16'h29b1, 16'h29ae, 16'h29ab, 16'h29a8, 16'h29a5, 16'h29a2, 16'h299f, 16'h299c, 16'h2999, 16'h2996, 16'h2993, 16'h2990, 16'h298d, 16'h298a, 16'h2987, 16'h2984, 16'h2981, 16'h297e, 16'h297b, 16'h2978, 16'h2975, 16'h2972, 16'h296f, 16'h296c, 16'h2969, 16'h2966, 16'h2963, 16'h2960, 16'h295d, 16'h295a, 16'h2957, 16'h2954, 16'h2951, 16'h294e, 16'h294b, 16'h2948, 16'h2945, 16'h2942, 16'h293f, 16'h293c, 16'h2939, 16'h2936, 16'h2933, 16'h2930, 16'h292d, 16'h292a, 16'h2927, 16'h2924, 16'h2921, 16'h291e, 16'h291b, 16'h2918, 16'h2915, 16'h2912, 16'h290f},
                                {16'h290c, 16'h2909, 16'h2906, 16'h2903, 16'h2900, 16'h28fd, 16'h28fa, 16'h28f7, 16'h28f4, 16'h28f1, 16'h28ee, 16'h28eb, 16'h28e8, 16'h28e5, 16'h28e2, 16'h28df, 16'h28dc, 16'h28d9, 16'h28d6, 16'h28d3, 16'h28d0, 16'h28cd, 16'h28ca, 16'h28c7, 16'h28c4, 16'h28c1, 16'h28be, 16'h28bb, 16'h28b8, 16'h28b5, 16'h28b2, 16'h28af, 16'h28ac, 16'h28a9, 16'h28a6, 16'h28a3, 16'h28a0, 16'h289d, 16'h289a, 16'h2897, 16'h2894, 16'h2891, 16'h288e, 16'h288b, 16'h2888, 16'h2885, 16'h2882, 16'h287f, 16'h287c, 16'h2879, 16'h2876, 16'h2873, 16'h2870, 16'h286d, 16'h286a, 16'h2867, 16'h2864, 16'h2861, 16'h285e, 16'h285b, 16'h2858, 16'h2855, 16'h2852, 16'h284f},
                                {16'h284c, 16'h2849, 16'h2846, 16'h2843, 16'h2840, 16'h283d, 16'h283a, 16'h2837, 16'h2834, 16'h2831, 16'h282e, 16'h282b, 16'h2828, 16'h2825, 16'h2822, 16'h281f, 16'h281c, 16'h2819, 16'h2816, 16'h2813, 16'h2810, 16'h280d, 16'h280a, 16'h2807, 16'h2804, 16'h2801, 16'h27fe, 16'h27fb, 16'h27f8, 16'h27f5, 16'h27f2, 16'h27ef, 16'h27ec, 16'h27e9, 16'h27e6, 16'h27e3, 16'h27e0, 16'h27dd, 16'h27da, 16'h27d7, 16'h27d4, 16'h27d1, 16'h27ce, 16'h27cb, 16'h27c8, 16'h27c5, 16'h27c2, 16'h27bf, 16'h27bc, 16'h27b9, 16'h27b6, 16'h27b3, 16'h27b0, 16'h27ad, 16'h27aa, 16'h27a7, 16'h27a4, 16'h27a1, 16'h279e, 16'h279b, 16'h2798, 16'h2795, 16'h2792, 16'h278f},
                                {16'h278c, 16'h2789, 16'h2786, 16'h2783, 16'h2780, 16'h277d, 16'h277a, 16'h2777, 16'h2774, 16'h2771, 16'h276e, 16'h276b, 16'h2768, 16'h2765, 16'h2762, 16'h275f, 16'h275c, 16'h2759, 16'h2756, 16'h2753, 16'h2750, 16'h274d, 16'h274a, 16'h2747, 16'h2744, 16'h2741, 16'h273e, 16'h273b, 16'h2738, 16'h2735, 16'h2732, 16'h272f, 16'h272c, 16'h2729, 16'h2726, 16'h2723, 16'h2720, 16'h271d, 16'h271a, 16'h2717, 16'h2714, 16'h2711, 16'h270e, 16'h270b, 16'h2708, 16'h2705, 16'h2702, 16'h26ff, 16'h26fc, 16'h26f9, 16'h26f6, 16'h26f3, 16'h26f0, 16'h26ed, 16'h26ea, 16'h26e7, 16'h26e4, 16'h26e1, 16'h26de, 16'h26db, 16'h26d8, 16'h26d5, 16'h26d2, 16'h26cf},
                                {16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc},
                                {16'h26cc, 16'h26cc, 16'h26cc, 16'h26cc, 16'h26c8, 16'h26c4, 16'h26c0, 16'h26bc, 16'h26b8, 16'h26b4, 16'h26b0, 16'h26ac, 16'h26a8, 16'h26a4, 16'h26a0, 16'h269c, 16'h2698, 16'h2694, 16'h2690, 16'h268c, 16'h2688, 16'h2684, 16'h2680, 16'h267c, 16'h2678, 16'h2674, 16'h2670, 16'h266c, 16'h2668, 16'h2664, 16'h2660, 16'h265c, 16'h2658, 16'h2654, 16'h2650, 16'h264c, 16'h2648, 16'h2644, 16'h2640, 16'h263c, 16'h2638, 16'h2634, 16'h2630, 16'h262c, 16'h2628, 16'h2624, 16'h2620, 16'h261c, 16'h2618, 16'h2614, 16'h2610, 16'h260c, 16'h2608, 16'h2604, 16'h2600, 16'h25fc, 16'h25f8, 16'h25f4, 16'h25f0, 16'h25ec, 16'h25e8, 16'h25e4, 16'h25e0, 16'h25dc},
                                {16'h25d8, 16'h25d4, 16'h25d0, 16'h25cc, 16'h25c8, 16'h25c4, 16'h25c0, 16'h25bc, 16'h25b8, 16'h25b4, 16'h25b0, 16'h25ac, 16'h25a8, 16'h25a4, 16'h25a0, 16'h259c, 16'h2598, 16'h2594, 16'h2590, 16'h258c, 16'h2588, 16'h2584, 16'h2580, 16'h257c, 16'h2578, 16'h2574, 16'h2570, 16'h256c, 16'h2568, 16'h2564, 16'h2560, 16'h255c, 16'h2558, 16'h2554, 16'h2550, 16'h254c, 16'h2548, 16'h2544, 16'h2540, 16'h253c, 16'h2538, 16'h2534, 16'h2530, 16'h252c, 16'h2528, 16'h2524, 16'h2520, 16'h251c, 16'h2518, 16'h2514, 16'h2510, 16'h250c, 16'h2508, 16'h2504, 16'h2500, 16'h24fc, 16'h24f8, 16'h24f4, 16'h24f0, 16'h24ec, 16'h24e8, 16'h24e4, 16'h24e0, 16'h24dc},
                                {16'h24d8, 16'h24d4, 16'h24d0, 16'h24cc, 16'h24c8, 16'h24c4, 16'h24c0, 16'h24bc, 16'h24b8, 16'h24b4, 16'h24b0, 16'h24ac, 16'h24a8, 16'h24a4, 16'h24a0, 16'h249c, 16'h2498, 16'h2494, 16'h2490, 16'h248c, 16'h2488, 16'h2484, 16'h2480, 16'h247c, 16'h2478, 16'h2474, 16'h2470, 16'h246c, 16'h2468, 16'h2464, 16'h2460, 16'h245c, 16'h2458, 16'h2454, 16'h2450, 16'h244c, 16'h2448, 16'h2444, 16'h2440, 16'h243c, 16'h2438, 16'h2434, 16'h2430, 16'h242c, 16'h2428, 16'h2424, 16'h2420, 16'h241c, 16'h2418, 16'h2414, 16'h2410, 16'h240c, 16'h2408, 16'h2404, 16'h2400, 16'h23fc, 16'h23f8, 16'h23f4, 16'h23f0, 16'h23ec, 16'h23e8, 16'h23e4, 16'h23e0, 16'h23dc},
                                {16'h23d8, 16'h23d4, 16'h23d0, 16'h23cc, 16'h23c8, 16'h23c4, 16'h23c0, 16'h23bc, 16'h23b8, 16'h23b4, 16'h23b0, 16'h23ac, 16'h23a8, 16'h23a4, 16'h23a0, 16'h239c, 16'h2398, 16'h2394, 16'h2390, 16'h238c, 16'h2388, 16'h2384, 16'h2380, 16'h237c, 16'h2378, 16'h2374, 16'h2370, 16'h236c, 16'h2368, 16'h2364, 16'h2360, 16'h235c, 16'h2358, 16'h2354, 16'h2350, 16'h234c, 16'h2348, 16'h2344, 16'h2340, 16'h233c, 16'h2338, 16'h2334, 16'h2330, 16'h232c, 16'h2328, 16'h2324, 16'h2320, 16'h231c, 16'h2318, 16'h2314, 16'h2310, 16'h230c, 16'h2308, 16'h2304, 16'h2300, 16'h22fc, 16'h22f8, 16'h22f4, 16'h22f0, 16'h22ec, 16'h22e8, 16'h22e4, 16'h22e0, 16'h22dc},
                                {16'h22d8, 16'h22d4, 16'h22d0, 16'h22cc, 16'h22c8, 16'h22c4, 16'h22c0, 16'h22bc, 16'h22b8, 16'h22b4, 16'h22b0, 16'h22ac, 16'h22a8, 16'h22a4, 16'h22a0, 16'h229c, 16'h2298, 16'h2294, 16'h2290, 16'h228c, 16'h2288, 16'h2284, 16'h2280, 16'h227c, 16'h2278, 16'h2274, 16'h2270, 16'h226c, 16'h2268, 16'h2264, 16'h2260, 16'h225c, 16'h2258, 16'h2254, 16'h2250, 16'h224c, 16'h2248, 16'h2244, 16'h2240, 16'h223c, 16'h2238, 16'h2234, 16'h2230, 16'h222c, 16'h2228, 16'h2224, 16'h2220, 16'h221c, 16'h2218, 16'h2214, 16'h2210, 16'h220c, 16'h2208, 16'h2204, 16'h2200, 16'h21fc, 16'h21f8, 16'h21f4, 16'h21f0, 16'h21ec, 16'h21e8, 16'h21e4, 16'h21e0, 16'h21dc},
                                {16'h21d8, 16'h21d4, 16'h21d0, 16'h21cc, 16'h21c8, 16'h21c4, 16'h21c0, 16'h21bc, 16'h21b8, 16'h21b4, 16'h21b0, 16'h21ac, 16'h21a8, 16'h21a4, 16'h21a0, 16'h219c, 16'h2198, 16'h2194, 16'h2190, 16'h218c, 16'h2188, 16'h2184, 16'h2180, 16'h217c, 16'h2178, 16'h2174, 16'h2170, 16'h216c, 16'h2168, 16'h2164, 16'h2160, 16'h215c, 16'h2158, 16'h2154, 16'h2150, 16'h214c, 16'h2148, 16'h2144, 16'h2140, 16'h213c, 16'h2138, 16'h2134, 16'h2130, 16'h212c, 16'h2128, 16'h2124, 16'h2120, 16'h211c, 16'h2118, 16'h2114, 16'h2110, 16'h210c, 16'h2108, 16'h2104, 16'h2100, 16'h20fc, 16'h20f8, 16'h20f4, 16'h20f0, 16'h20ec, 16'h20e8, 16'h20e4, 16'h20e0, 16'h20dc},
                                {16'h20d8, 16'h20d4, 16'h20d0, 16'h20cc, 16'h20c8, 16'h20c4, 16'h20c0, 16'h20bc, 16'h20b8, 16'h20b4, 16'h20b0, 16'h20ac, 16'h20a8, 16'h20a4, 16'h20a0, 16'h209c, 16'h2098, 16'h2094, 16'h2090, 16'h208c, 16'h2088, 16'h2084, 16'h2080, 16'h207c, 16'h2078, 16'h2074, 16'h2070, 16'h206c, 16'h2068, 16'h2064, 16'h2060, 16'h205c, 16'h2058, 16'h2054, 16'h2050, 16'h204c, 16'h2048, 16'h2044, 16'h2040, 16'h203c, 16'h2038, 16'h2034, 16'h2030, 16'h202c, 16'h2028, 16'h2024, 16'h2020, 16'h201c, 16'h2018, 16'h2014, 16'h2010, 16'h200c, 16'h2008, 16'h2004, 16'h2000, 16'h1ffc, 16'h1ff8, 16'h1ff4, 16'h1ff0, 16'h1fec, 16'h1fe8, 16'h1fe4, 16'h1fe0, 16'h1fdc},
                                {16'h1fd8, 16'h1fd4, 16'h1fd0, 16'h1fcc, 16'h1fc8, 16'h1fc4, 16'h1fc0, 16'h1fbc, 16'h1fb8, 16'h1fb4, 16'h1fb0, 16'h1fac, 16'h1fa8, 16'h1fa4, 16'h1fa0, 16'h1f9c, 16'h1f98, 16'h1f94, 16'h1f90, 16'h1f8c, 16'h1f88, 16'h1f84, 16'h1f80, 16'h1f7c, 16'h1f78, 16'h1f74, 16'h1f70, 16'h1f6c, 16'h1f68, 16'h1f64, 16'h1f60, 16'h1f5c, 16'h1f58, 16'h1f54, 16'h1f50, 16'h1f4c, 16'h1f48, 16'h1f44, 16'h1f40, 16'h1f3c, 16'h1f38, 16'h1f34, 16'h1f30, 16'h1f2c, 16'h1f28, 16'h1f24, 16'h1f20, 16'h1f1c, 16'h1f18, 16'h1f14, 16'h1f10, 16'h1f0c, 16'h1f08, 16'h1f04, 16'h1f00, 16'h1efc, 16'h1ef8, 16'h1ef4, 16'h1ef0, 16'h1eec, 16'h1ee8, 16'h1ee4, 16'h1ee0, 16'h1edc},
                                {16'h1ed8, 16'h1ed4, 16'h1ed0, 16'h1ecc, 16'h1ec8, 16'h1ec4, 16'h1ec0, 16'h1ebc, 16'h1eb8, 16'h1eb4, 16'h1eb0, 16'h1eac, 16'h1ea8, 16'h1ea4, 16'h1ea0, 16'h1e9c, 16'h1e98, 16'h1e94, 16'h1e90, 16'h1e8c, 16'h1e88, 16'h1e84, 16'h1e80, 16'h1e7c, 16'h1e78, 16'h1e74, 16'h1e70, 16'h1e6c, 16'h1e68, 16'h1e64, 16'h1e60, 16'h1e5c, 16'h1e58, 16'h1e54, 16'h1e50, 16'h1e4c, 16'h1e48, 16'h1e44, 16'h1e40, 16'h1e3c, 16'h1e38, 16'h1e34, 16'h1e30, 16'h1e2c, 16'h1e28, 16'h1e24, 16'h1e20, 16'h1e1c, 16'h1e18, 16'h1e14, 16'h1e10, 16'h1e0c, 16'h1e08, 16'h1e04, 16'h1e00, 16'h1dfc, 16'h1df8, 16'h1df4, 16'h1df0, 16'h1dec, 16'h1de8, 16'h1de4, 16'h1de0, 16'h1ddc},
                                {16'h1dd8, 16'h1dd4, 16'h1dd0, 16'h1dcc, 16'h1dc8, 16'h1dc4, 16'h1dc0, 16'h1dbc, 16'h1db8, 16'h1db4, 16'h1db0, 16'h1dac, 16'h1da8, 16'h1da4, 16'h1da0, 16'h1d9c, 16'h1d98, 16'h1d94, 16'h1d90, 16'h1d8c, 16'h1d88, 16'h1d84, 16'h1d80, 16'h1d7c, 16'h1d78, 16'h1d74, 16'h1d70, 16'h1d6c, 16'h1d68, 16'h1d64, 16'h1d60, 16'h1d5c, 16'h1d58, 16'h1d54, 16'h1d50, 16'h1d4c, 16'h1d48, 16'h1d44, 16'h1d40, 16'h1d3c, 16'h1d38, 16'h1d34, 16'h1d30, 16'h1d2c, 16'h1d28, 16'h1d24, 16'h1d20, 16'h1d1c, 16'h1d18, 16'h1d14, 16'h1d10, 16'h1d0c, 16'h1d08, 16'h1d04, 16'h1d00, 16'h1cfc, 16'h1cf8, 16'h1cf4, 16'h1cf0, 16'h1cec, 16'h1ce8, 16'h1ce4, 16'h1ce0, 16'h1cdc},
                                {16'h1cd8, 16'h1cd4, 16'h1cd0, 16'h1ccc, 16'h1cc8, 16'h1cc4, 16'h1cc0, 16'h1cbc, 16'h1cb8, 16'h1cb4, 16'h1cb0, 16'h1cac, 16'h1ca8, 16'h1ca4, 16'h1ca0, 16'h1c9c, 16'h1c98, 16'h1c94, 16'h1c90, 16'h1c8c, 16'h1c88, 16'h1c84, 16'h1c80, 16'h1c7c, 16'h1c78, 16'h1c74, 16'h1c70, 16'h1c6c, 16'h1c68, 16'h1c64, 16'h1c60, 16'h1c5c, 16'h1c58, 16'h1c54, 16'h1c50, 16'h1c4c, 16'h1c48, 16'h1c44, 16'h1c40, 16'h1c3c, 16'h1c38, 16'h1c34, 16'h1c30, 16'h1c2c, 16'h1c28, 16'h1c24, 16'h1c20, 16'h1c1c, 16'h1c18, 16'h1c14, 16'h1c10, 16'h1c0c, 16'h1c08, 16'h1c04, 16'h1c00, 16'h1bfc, 16'h1bf8, 16'h1bf4, 16'h1bf0, 16'h1bec, 16'h1be8, 16'h1be4, 16'h1be0, 16'h1bdc},
                                {16'h1bd8, 16'h1bd4, 16'h1bd0, 16'h1bcc, 16'h1bc8, 16'h1bc4, 16'h1bc0, 16'h1bbc, 16'h1bb8, 16'h1bb4, 16'h1bb0, 16'h1bac, 16'h1ba8, 16'h1ba4, 16'h1ba0, 16'h1b9c, 16'h1b98, 16'h1b94, 16'h1b90, 16'h1b8c, 16'h1b88, 16'h1b84, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80},
                                {16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b80, 16'h1b7e, 16'h1b7b, 16'h1b78, 16'h1b75, 16'h1b72},
                                {16'h1b6f, 16'h1b6c, 16'h1b69, 16'h1b66, 16'h1b63, 16'h1b60, 16'h1b5d, 16'h1b5a, 16'h1b57, 16'h1b54, 16'h1b51, 16'h1b4e, 16'h1b4b, 16'h1b48, 16'h1b45, 16'h1b42, 16'h1b3f, 16'h1b3c, 16'h1b39, 16'h1b36, 16'h1b33, 16'h1b30, 16'h1b2d, 16'h1b2a, 16'h1b27, 16'h1b24, 16'h1b21, 16'h1b1e, 16'h1b1b, 16'h1b18, 16'h1b15, 16'h1b12, 16'h1b0f, 16'h1b0c, 16'h1b09, 16'h1b06, 16'h1b03, 16'h1b00, 16'h1afd, 16'h1afa, 16'h1af7, 16'h1af4, 16'h1af1, 16'h1aee, 16'h1aeb, 16'h1ae8, 16'h1ae5, 16'h1ae2, 16'h1adf, 16'h1adc, 16'h1ad9, 16'h1ad6, 16'h1ad3, 16'h1ad0, 16'h1acd, 16'h1aca, 16'h1ac7, 16'h1ac4, 16'h1ac1, 16'h1abe, 16'h1abb, 16'h1ab8, 16'h1ab5, 16'h1ab2},
                                {16'h1aaf, 16'h1aac, 16'h1aa9, 16'h1aa6, 16'h1aa3, 16'h1aa0, 16'h1a9d, 16'h1a9a, 16'h1a97, 16'h1a94, 16'h1a91, 16'h1a8e, 16'h1a8b, 16'h1a88, 16'h1a85, 16'h1a82, 16'h1a7f, 16'h1a7c, 16'h1a79, 16'h1a76, 16'h1a73, 16'h1a70, 16'h1a6d, 16'h1a6a, 16'h1a67, 16'h1a64, 16'h1a61, 16'h1a5e, 16'h1a5b, 16'h1a58, 16'h1a55, 16'h1a52, 16'h1a4f, 16'h1a4c, 16'h1a49, 16'h1a46, 16'h1a43, 16'h1a40, 16'h1a3d, 16'h1a3a, 16'h1a37, 16'h1a34, 16'h1a31, 16'h1a2e, 16'h1a2b, 16'h1a28, 16'h1a25, 16'h1a22, 16'h1a1f, 16'h1a1c, 16'h1a19, 16'h1a16, 16'h1a13, 16'h1a10, 16'h1a0d, 16'h1a0a, 16'h1a07, 16'h1a04, 16'h1a01, 16'h19fe, 16'h19fb, 16'h19f8, 16'h19f5, 16'h19f2},
                                {16'h19ef, 16'h19ec, 16'h19e9, 16'h19e6, 16'h19e3, 16'h19e0, 16'h19dd, 16'h19da, 16'h19d7, 16'h19d4, 16'h19d1, 16'h19ce, 16'h19cb, 16'h19c8, 16'h19c5, 16'h19c2, 16'h19bf, 16'h19bc, 16'h19b9, 16'h19b6, 16'h19b3, 16'h19b0, 16'h19ad, 16'h19aa, 16'h19a7, 16'h19a4, 16'h19a1, 16'h199e, 16'h199b, 16'h1998, 16'h1995, 16'h1992, 16'h198f, 16'h198c, 16'h1989, 16'h1986, 16'h1983, 16'h1980, 16'h197d, 16'h197a, 16'h1977, 16'h1974, 16'h1971, 16'h196e, 16'h196b, 16'h1968, 16'h1965, 16'h1962, 16'h195f, 16'h195c, 16'h1959, 16'h1956, 16'h1953, 16'h1950, 16'h194d, 16'h194a, 16'h1947, 16'h1944, 16'h1941, 16'h193e, 16'h193b, 16'h1938, 16'h1935, 16'h1932},
                                {16'h192f, 16'h192c, 16'h1929, 16'h1926, 16'h1923, 16'h1920, 16'h191d, 16'h191a, 16'h1917, 16'h1914, 16'h1911, 16'h190e, 16'h190b, 16'h1908, 16'h1905, 16'h1902, 16'h18ff, 16'h18fc, 16'h18f9, 16'h18f6, 16'h18f3, 16'h18f0, 16'h18ed, 16'h18ea, 16'h18e7, 16'h18e4, 16'h18e1, 16'h18de, 16'h18db, 16'h18d8, 16'h18d5, 16'h18d2, 16'h18cf, 16'h18cc, 16'h18c9, 16'h18c6, 16'h18c3, 16'h18c0, 16'h18bd, 16'h18ba, 16'h18b7, 16'h18b4, 16'h18b1, 16'h18ae, 16'h18ab, 16'h18a8, 16'h18a5, 16'h18a2, 16'h189f, 16'h189c, 16'h1899, 16'h1896, 16'h1893, 16'h1890, 16'h188d, 16'h188a, 16'h1887, 16'h1884, 16'h1881, 16'h187e, 16'h187b, 16'h1878, 16'h1875, 16'h1872},
                                {16'h186f, 16'h186c, 16'h1869, 16'h1866, 16'h1863, 16'h1860, 16'h185d, 16'h185a, 16'h1857, 16'h1854, 16'h1851, 16'h184e, 16'h184b, 16'h1848, 16'h1845, 16'h1842, 16'h183f, 16'h183c, 16'h1839, 16'h1836, 16'h1833, 16'h1830, 16'h182d, 16'h182a, 16'h1827, 16'h1824, 16'h1821, 16'h181e, 16'h181b, 16'h1818, 16'h1815, 16'h1812, 16'h180f, 16'h180c, 16'h1809, 16'h1806, 16'h1803, 16'h1800, 16'h17fd, 16'h17fa, 16'h17f7, 16'h17f4, 16'h17f1, 16'h17ee, 16'h17eb, 16'h17e8, 16'h17e5, 16'h17e2, 16'h17df, 16'h17dc, 16'h17d9, 16'h17d6, 16'h17d3, 16'h17d0, 16'h17cd, 16'h17ca, 16'h17c7, 16'h17c4, 16'h17c1, 16'h17be, 16'h17bb, 16'h17b8, 16'h17b5, 16'h17b2},
                                {16'h17af, 16'h17ac, 16'h17a9, 16'h17a6, 16'h17a3, 16'h17a0, 16'h179d, 16'h179a, 16'h1797, 16'h1794, 16'h1791, 16'h178e, 16'h178b, 16'h1788, 16'h1785, 16'h1782, 16'h177f, 16'h177c, 16'h1779, 16'h1776, 16'h1773, 16'h1770, 16'h176d, 16'h176a, 16'h1767, 16'h1764, 16'h1761, 16'h175e, 16'h175b, 16'h1758, 16'h1755, 16'h1752, 16'h174f, 16'h174c, 16'h1749, 16'h1746, 16'h1743, 16'h1740, 16'h173d, 16'h173a, 16'h1737, 16'h1734, 16'h1731, 16'h172e, 16'h172b, 16'h1728, 16'h1725, 16'h1722, 16'h171f, 16'h171c, 16'h1719, 16'h1716, 16'h1713, 16'h1710, 16'h170d, 16'h170a, 16'h1707, 16'h1704, 16'h1701, 16'h16fe, 16'h16fb, 16'h16f8, 16'h16f5, 16'h16f2},
                                {16'h16ef, 16'h16ec, 16'h16e9, 16'h16e6, 16'h16e3, 16'h16e0, 16'h16dd, 16'h16da, 16'h16d7, 16'h16d4, 16'h16d1, 16'h16ce, 16'h16cb, 16'h16c8, 16'h16c5, 16'h16c2, 16'h16bf, 16'h16bc, 16'h16b9, 16'h16b6, 16'h16b3, 16'h16b0, 16'h16ad, 16'h16aa, 16'h16a7, 16'h16a4, 16'h16a1, 16'h169e, 16'h169b, 16'h1698, 16'h1695, 16'h1692, 16'h168f, 16'h168c, 16'h1689, 16'h1686, 16'h1683, 16'h1680, 16'h167d, 16'h167a, 16'h1677, 16'h1674, 16'h1671, 16'h166e, 16'h166b, 16'h1668, 16'h1665, 16'h1662, 16'h165f, 16'h165c, 16'h1659, 16'h1656, 16'h1653, 16'h1650, 16'h164d, 16'h164a, 16'h1647, 16'h1644, 16'h1641, 16'h163e, 16'h163b, 16'h1638, 16'h1635, 16'h1632},
                                {16'h162f, 16'h162c, 16'h1629, 16'h1626, 16'h1623, 16'h1620, 16'h161d, 16'h161a, 16'h1617, 16'h1614, 16'h1611, 16'h160e, 16'h160b, 16'h1608, 16'h1605, 16'h1602, 16'h15ff, 16'h15fc, 16'h15f9, 16'h15f6, 16'h15f3, 16'h15f0, 16'h15ed, 16'h15ea, 16'h15e7, 16'h15e4, 16'h15e1, 16'h15de, 16'h15db, 16'h15d8, 16'h15d5, 16'h15d2, 16'h15cf, 16'h15cc, 16'h15c9, 16'h15c6, 16'h15c3, 16'h15c0, 16'h15bd, 16'h15ba, 16'h15b7, 16'h15b4, 16'h15b1, 16'h15ae, 16'h15ab, 16'h15a8, 16'h15a5, 16'h15a2, 16'h159f, 16'h159c, 16'h1599, 16'h1596, 16'h1593, 16'h1590, 16'h158d, 16'h158a, 16'h1587, 16'h1584, 16'h1581, 16'h157e, 16'h157b, 16'h1578, 16'h1575, 16'h1572},
                                {16'h156f, 16'h156c, 16'h1569, 16'h1566, 16'h1563, 16'h1560, 16'h155d, 16'h155a, 16'h1557, 16'h1554, 16'h1551, 16'h154e, 16'h154b, 16'h1548, 16'h1545, 16'h1542, 16'h153f, 16'h153c, 16'h1539, 16'h1536, 16'h1533, 16'h1530, 16'h152d, 16'h152a, 16'h1527, 16'h1524, 16'h1521, 16'h151e, 16'h151b, 16'h1518, 16'h1515, 16'h1512, 16'h150f, 16'h150c, 16'h1509, 16'h1506, 16'h1503, 16'h1500, 16'h14fd, 16'h14fa, 16'h14f7, 16'h14f4, 16'h14f1, 16'h14ee, 16'h14eb, 16'h14e8, 16'h14e5, 16'h14e2, 16'h14df, 16'h14dc, 16'h14d9, 16'h14d6, 16'h14d3, 16'h14d0, 16'h14cd, 16'h14ca, 16'h14c7, 16'h14c4, 16'h14c1, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be},
                                {16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be},
                                {16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14be, 16'h14bb, 16'h14b8, 16'h14b5, 16'h14b2, 16'h14af, 16'h14ac, 16'h14a9, 16'h14a6, 16'h14a3, 16'h14a0, 16'h149d, 16'h149a, 16'h1497, 16'h1494, 16'h1491, 16'h148e, 16'h148b, 16'h1488, 16'h1485, 16'h1482, 16'h147f, 16'h147c, 16'h1479, 16'h1476, 16'h1473, 16'h1470, 16'h146d, 16'h146a, 16'h1467, 16'h1464, 16'h1461, 16'h145e},
                                {16'h145b, 16'h1458, 16'h1455, 16'h1452, 16'h144f, 16'h144c, 16'h1449, 16'h1446, 16'h1443, 16'h1440, 16'h143d, 16'h143a, 16'h1437, 16'h1434, 16'h1431, 16'h142e, 16'h142b, 16'h1428, 16'h1425, 16'h1422, 16'h141f, 16'h141c, 16'h1419, 16'h1416, 16'h1413, 16'h1410, 16'h140d, 16'h140a, 16'h1407, 16'h1404, 16'h1401, 16'h13fe, 16'h13fb, 16'h13f8, 16'h13f5, 16'h13f2, 16'h13ef, 16'h13ec, 16'h13e9, 16'h13e6, 16'h13e3, 16'h13e0, 16'h13dd, 16'h13da, 16'h13d7, 16'h13d4, 16'h13d1, 16'h13ce, 16'h13cb, 16'h13c8, 16'h13c5, 16'h13c2, 16'h13bf, 16'h13bc, 16'h13b9, 16'h13b6, 16'h13b3, 16'h13b0, 16'h13ad, 16'h13aa, 16'h13a7, 16'h13a4, 16'h13a1, 16'h139e},
                                {16'h139b, 16'h1398, 16'h1395, 16'h1392, 16'h138f, 16'h138c, 16'h1389, 16'h1386, 16'h1383, 16'h1380, 16'h137d, 16'h137a, 16'h1377, 16'h1374, 16'h1371, 16'h136e, 16'h136b, 16'h1368, 16'h1365, 16'h1362, 16'h135f, 16'h135c, 16'h1359, 16'h1356, 16'h1353, 16'h1350, 16'h134d, 16'h134a, 16'h1347, 16'h1344, 16'h1341, 16'h133e, 16'h133b, 16'h1338, 16'h1335, 16'h1332, 16'h132f, 16'h132c, 16'h1329, 16'h1326, 16'h1323, 16'h1320, 16'h131d, 16'h131a, 16'h1317, 16'h1314, 16'h1311, 16'h130e, 16'h130b, 16'h1308, 16'h1305, 16'h1302, 16'h12ff, 16'h12fc, 16'h12f9, 16'h12f6, 16'h12f3, 16'h12f0, 16'h12ed, 16'h12ea, 16'h12e7, 16'h12e4, 16'h12e1, 16'h12de},
                                {16'h12db, 16'h12d8, 16'h12d5, 16'h12d2, 16'h12cf, 16'h12cc, 16'h12c9, 16'h12c6, 16'h12c3, 16'h12c0, 16'h12bd, 16'h12ba, 16'h12b7, 16'h12b4, 16'h12b1, 16'h12ae, 16'h12ab, 16'h12a8, 16'h12a5, 16'h12a2, 16'h129f, 16'h129c, 16'h1299, 16'h1296, 16'h1293, 16'h1290, 16'h128d, 16'h128a, 16'h1287, 16'h1284, 16'h1281, 16'h127e, 16'h127b, 16'h1278, 16'h1275, 16'h1272, 16'h126f, 16'h126c, 16'h1269, 16'h1266, 16'h1263, 16'h1260, 16'h125d, 16'h125a, 16'h1257, 16'h1254, 16'h1251, 16'h124e, 16'h124b, 16'h1248, 16'h1245, 16'h1242, 16'h123f, 16'h123c, 16'h1239, 16'h1236, 16'h1233, 16'h1230, 16'h122d, 16'h122a, 16'h1227, 16'h1224, 16'h1221, 16'h121e},
                                {16'h121b, 16'h1218, 16'h1215, 16'h1212, 16'h120f, 16'h120c, 16'h1209, 16'h1206, 16'h1203, 16'h1200, 16'h11fd, 16'h11fa, 16'h11f7, 16'h11f4, 16'h11f1, 16'h11ee, 16'h11eb, 16'h11e8, 16'h11e5, 16'h11e2, 16'h11df, 16'h11dc, 16'h11d9, 16'h11d6, 16'h11d3, 16'h11d0, 16'h11cd, 16'h11ca, 16'h11c7, 16'h11c4, 16'h11c1, 16'h11be, 16'h11bb, 16'h11b8, 16'h11b5, 16'h11b2, 16'h11af, 16'h11ac, 16'h11a9, 16'h11a6, 16'h11a3, 16'h11a0, 16'h119d, 16'h119a, 16'h1197, 16'h1194, 16'h1191, 16'h118e, 16'h118b, 16'h1188, 16'h1185, 16'h1182, 16'h117f, 16'h117c, 16'h1179, 16'h1176, 16'h1173, 16'h1170, 16'h116d, 16'h116a, 16'h1167, 16'h1164, 16'h1161, 16'h115e},
                                {16'h115b, 16'h1158, 16'h1155, 16'h1152, 16'h114f, 16'h114c, 16'h1149, 16'h1146, 16'h1143, 16'h1140, 16'h113d, 16'h113a, 16'h1137, 16'h1134, 16'h1131, 16'h112e, 16'h112b, 16'h1128, 16'h1125, 16'h1122, 16'h111f, 16'h111c, 16'h1119, 16'h1116, 16'h1113, 16'h1110, 16'h110d, 16'h110a, 16'h1107, 16'h1104, 16'h1101, 16'h10fe, 16'h10fb, 16'h10f8, 16'h10f5, 16'h10f2, 16'h10ef, 16'h10ec, 16'h10e9, 16'h10e6, 16'h10e3, 16'h10e0, 16'h10dd, 16'h10da, 16'h10d7, 16'h10d4, 16'h10d1, 16'h10ce, 16'h10cb, 16'h10c8, 16'h10c5, 16'h10c2, 16'h10bf, 16'h10bc, 16'h10b9, 16'h10b6, 16'h10b3, 16'h10b0, 16'h10ad, 16'h10aa, 16'h10a7, 16'h10a4, 16'h10a1, 16'h109e},
                                {16'h109b, 16'h1098, 16'h1095, 16'h1092, 16'h108f, 16'h108c, 16'h1089, 16'h1086, 16'h1083, 16'h1080, 16'h107d, 16'h107a, 16'h1077, 16'h1074, 16'h1071, 16'h106e, 16'h106b, 16'h1068, 16'h1065, 16'h1062, 16'h105f, 16'h105c, 16'h1059, 16'h1056, 16'h1053, 16'h1050, 16'h104d, 16'h104a, 16'h1047, 16'h1044, 16'h1041, 16'h103e, 16'h103b, 16'h1038, 16'h1035, 16'h1032, 16'h102f, 16'h102c, 16'h1029, 16'h1026, 16'h1023, 16'h1020, 16'h101d, 16'h101a, 16'h1017, 16'h1014, 16'h1011, 16'h100e, 16'h100b, 16'h1008, 16'h1005, 16'h1002, 16'h0fff, 16'h0ffc, 16'h0ff9, 16'h0ff6, 16'h0ff3, 16'h0ff0, 16'h0fed, 16'h0fea, 16'h0fe7, 16'h0fe4, 16'h0fe1, 16'h0fde},
                                {16'h0fdb, 16'h0fd8, 16'h0fd5, 16'h0fd2, 16'h0fcf, 16'h0fcc, 16'h0fc9, 16'h0fc6, 16'h0fc3, 16'h0fc0, 16'h0fbd, 16'h0fba, 16'h0fb7, 16'h0fb4, 16'h0fb1, 16'h0fae, 16'h0fab, 16'h0fa8, 16'h0fa5, 16'h0fa2, 16'h0f9f, 16'h0f9c, 16'h0f99, 16'h0f96, 16'h0f93, 16'h0f90, 16'h0f8d, 16'h0f8a, 16'h0f87, 16'h0f84, 16'h0f81, 16'h0f7e, 16'h0f7b, 16'h0f78, 16'h0f75, 16'h0f72, 16'h0f6f, 16'h0f6c, 16'h0f69, 16'h0f66, 16'h0f63, 16'h0f60, 16'h0f5d, 16'h0f5a, 16'h0f57, 16'h0f54, 16'h0f51, 16'h0f4e, 16'h0f4b, 16'h0f48, 16'h0f45, 16'h0f42, 16'h0f3f, 16'h0f3c, 16'h0f39, 16'h0f36, 16'h0f33, 16'h0f30, 16'h0f2d, 16'h0f2a, 16'h0f27, 16'h0f24, 16'h0f21, 16'h0f1e},
                                {16'h0f1b, 16'h0f18, 16'h0f15, 16'h0f12, 16'h0f0f, 16'h0f0c, 16'h0f09, 16'h0f06, 16'h0f03, 16'h0f00, 16'h0efd, 16'h0efa, 16'h0ef7, 16'h0ef4, 16'h0ef1, 16'h0eee, 16'h0eeb, 16'h0ee8, 16'h0ee5, 16'h0ee2, 16'h0edf, 16'h0edc, 16'h0ed9, 16'h0ed6, 16'h0ed3, 16'h0ed0, 16'h0ecd, 16'h0eca, 16'h0ec7, 16'h0ec4, 16'h0ec1, 16'h0ebe, 16'h0ebb, 16'h0eb8, 16'h0eb5, 16'h0eb2, 16'h0eaf, 16'h0eac, 16'h0ea9, 16'h0ea6, 16'h0ea3, 16'h0ea0, 16'h0e9d, 16'h0e9a, 16'h0e97, 16'h0e94, 16'h0e91, 16'h0e8e, 16'h0e8b, 16'h0e88, 16'h0e85, 16'h0e82, 16'h0e7f, 16'h0e7c, 16'h0e79, 16'h0e76, 16'h0e73, 16'h0e70, 16'h0e6d, 16'h0e6a, 16'h0e67, 16'h0e64, 16'h0e61, 16'h0e5e},
                                {16'h0e5b, 16'h0e58, 16'h0e55, 16'h0e52, 16'h0e4f, 16'h0e4c, 16'h0e49, 16'h0e46, 16'h0e43, 16'h0e40, 16'h0e3d, 16'h0e3a, 16'h0e37, 16'h0e34, 16'h0e31, 16'h0e2e, 16'h0e2b, 16'h0e28, 16'h0e25, 16'h0e22, 16'h0e1f, 16'h0e1c, 16'h0e19, 16'h0e16, 16'h0e13, 16'h0e10, 16'h0e0d, 16'h0e0a, 16'h0e07, 16'h0e04, 16'h0e01, 16'h0dfe, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb},
                                {16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfb, 16'h0dfa, 16'h0df9, 16'h0df8, 16'h0df7, 16'h0df6, 16'h0df5, 16'h0df4, 16'h0df3, 16'h0df2, 16'h0df1, 16'h0df0, 16'h0def, 16'h0dee, 16'h0ded, 16'h0dec, 16'h0deb, 16'h0dea, 16'h0de9, 16'h0de8, 16'h0de7, 16'h0de6, 16'h0de5, 16'h0de4},
                                {16'h0de3, 16'h0de2, 16'h0de1, 16'h0de0, 16'h0ddf, 16'h0dde, 16'h0ddd, 16'h0ddc, 16'h0ddb, 16'h0dda, 16'h0dd9, 16'h0dd8, 16'h0dd7, 16'h0dd6, 16'h0dd5, 16'h0dd4, 16'h0dd3, 16'h0dd2, 16'h0dd1, 16'h0dd0, 16'h0dcf, 16'h0dce, 16'h0dcd, 16'h0dcc, 16'h0dcb, 16'h0dca, 16'h0dc9, 16'h0dc8, 16'h0dc7, 16'h0dc6, 16'h0dc5, 16'h0dc4, 16'h0dc3, 16'h0dc2, 16'h0dc1, 16'h0dc0, 16'h0dbf, 16'h0dbe, 16'h0dbd, 16'h0dbc, 16'h0dbb, 16'h0dba, 16'h0db9, 16'h0db8, 16'h0db7, 16'h0db6, 16'h0db5, 16'h0db4, 16'h0db3, 16'h0db2, 16'h0db1, 16'h0db0, 16'h0daf, 16'h0dae, 16'h0dad, 16'h0dac, 16'h0dab, 16'h0daa, 16'h0da9, 16'h0da8, 16'h0da7, 16'h0da6, 16'h0da5, 16'h0da4},
                                {16'h0da3, 16'h0da2, 16'h0da1, 16'h0da0, 16'h0d9f, 16'h0d9e, 16'h0d9d, 16'h0d9c, 16'h0d9b, 16'h0d9a, 16'h0d99, 16'h0d98, 16'h0d97, 16'h0d96, 16'h0d95, 16'h0d94, 16'h0d93, 16'h0d92, 16'h0d91, 16'h0d90, 16'h0d8f, 16'h0d8e, 16'h0d8d, 16'h0d8c, 16'h0d8b, 16'h0d8a, 16'h0d89, 16'h0d88, 16'h0d87, 16'h0d86, 16'h0d85, 16'h0d84, 16'h0d83, 16'h0d82, 16'h0d81, 16'h0d80, 16'h0d7f, 16'h0d7e, 16'h0d7d, 16'h0d7c, 16'h0d7b, 16'h0d7a, 16'h0d79, 16'h0d78, 16'h0d77, 16'h0d76, 16'h0d75, 16'h0d74, 16'h0d73, 16'h0d72, 16'h0d71, 16'h0d70, 16'h0d6f, 16'h0d6e, 16'h0d6d, 16'h0d6c, 16'h0d6b, 16'h0d6a, 16'h0d69, 16'h0d68, 16'h0d67, 16'h0d66, 16'h0d65, 16'h0d64},
                                {16'h0d63, 16'h0d62, 16'h0d61, 16'h0d60, 16'h0d5f, 16'h0d5e, 16'h0d5d, 16'h0d5c, 16'h0d5b, 16'h0d5a, 16'h0d59, 16'h0d58, 16'h0d57, 16'h0d56, 16'h0d55, 16'h0d54, 16'h0d53, 16'h0d52, 16'h0d51, 16'h0d50, 16'h0d4f, 16'h0d4e, 16'h0d4d, 16'h0d4c, 16'h0d4b, 16'h0d4a, 16'h0d49, 16'h0d48, 16'h0d47, 16'h0d46, 16'h0d45, 16'h0d44, 16'h0d43, 16'h0d42, 16'h0d41, 16'h0d40, 16'h0d3f, 16'h0d3e, 16'h0d3d, 16'h0d3c, 16'h0d3b, 16'h0d3a, 16'h0d39, 16'h0d38, 16'h0d37, 16'h0d36, 16'h0d35, 16'h0d34, 16'h0d33, 16'h0d32, 16'h0d31, 16'h0d30, 16'h0d2f, 16'h0d2e, 16'h0d2d, 16'h0d2c, 16'h0d2b, 16'h0d2a, 16'h0d29, 16'h0d28, 16'h0d27, 16'h0d26, 16'h0d25, 16'h0d24},
                                {16'h0d23, 16'h0d22, 16'h0d21, 16'h0d20, 16'h0d1f, 16'h0d1e, 16'h0d1d, 16'h0d1c, 16'h0d1b, 16'h0d1a, 16'h0d19, 16'h0d18, 16'h0d17, 16'h0d16, 16'h0d15, 16'h0d14, 16'h0d13, 16'h0d12, 16'h0d11, 16'h0d10, 16'h0d0f, 16'h0d0e, 16'h0d0d, 16'h0d0c, 16'h0d0b, 16'h0d0a, 16'h0d09, 16'h0d08, 16'h0d07, 16'h0d06, 16'h0d05, 16'h0d04, 16'h0d03, 16'h0d02, 16'h0d01, 16'h0d00, 16'h0cff, 16'h0cfe, 16'h0cfd, 16'h0cfc, 16'h0cfb, 16'h0cfa, 16'h0cf9, 16'h0cf8, 16'h0cf7, 16'h0cf6, 16'h0cf5, 16'h0cf4, 16'h0cf3, 16'h0cf2, 16'h0cf1, 16'h0cf0, 16'h0cef, 16'h0cee, 16'h0ced, 16'h0cec, 16'h0ceb, 16'h0cea, 16'h0ce9, 16'h0ce8, 16'h0ce7, 16'h0ce6, 16'h0ce5, 16'h0ce4},
                                {16'h0ce3, 16'h0ce2, 16'h0ce1, 16'h0ce0, 16'h0cdf, 16'h0cde, 16'h0cdd, 16'h0cdc, 16'h0cdb, 16'h0cda, 16'h0cd9, 16'h0cd8, 16'h0cd7, 16'h0cd6, 16'h0cd5, 16'h0cd4, 16'h0cd3, 16'h0cd2, 16'h0cd1, 16'h0cd0, 16'h0ccf, 16'h0cce, 16'h0ccd, 16'h0ccc, 16'h0ccb, 16'h0cca, 16'h0cc9, 16'h0cc8, 16'h0cc7, 16'h0cc6, 16'h0cc5, 16'h0cc4, 16'h0cc3, 16'h0cc2, 16'h0cc1, 16'h0cc0, 16'h0cbf, 16'h0cbe, 16'h0cbd, 16'h0cbc, 16'h0cbb, 16'h0cba, 16'h0cb9, 16'h0cb8, 16'h0cb7, 16'h0cb6, 16'h0cb5, 16'h0cb4, 16'h0cb3, 16'h0cb2, 16'h0cb1, 16'h0cb0, 16'h0caf, 16'h0cae, 16'h0cad, 16'h0cac, 16'h0cab, 16'h0caa, 16'h0ca9, 16'h0ca8, 16'h0ca7, 16'h0ca6, 16'h0ca5, 16'h0ca4},
                                {16'h0ca3, 16'h0ca2, 16'h0ca1, 16'h0ca0, 16'h0c9f, 16'h0c9e, 16'h0c9d, 16'h0c9c, 16'h0c9b, 16'h0c9a, 16'h0c99, 16'h0c98, 16'h0c97, 16'h0c96, 16'h0c95, 16'h0c94, 16'h0c93, 16'h0c92, 16'h0c91, 16'h0c90, 16'h0c8f, 16'h0c8e, 16'h0c8d, 16'h0c8c, 16'h0c8b, 16'h0c8a, 16'h0c89, 16'h0c88, 16'h0c87, 16'h0c86, 16'h0c85, 16'h0c84, 16'h0c83, 16'h0c82, 16'h0c81, 16'h0c80, 16'h0c7f, 16'h0c7e, 16'h0c7d, 16'h0c7c, 16'h0c7b, 16'h0c7a, 16'h0c79, 16'h0c78, 16'h0c77, 16'h0c76, 16'h0c75, 16'h0c74, 16'h0c73, 16'h0c72, 16'h0c71, 16'h0c70, 16'h0c6f, 16'h0c6e, 16'h0c6d, 16'h0c6c, 16'h0c6b, 16'h0c6a, 16'h0c69, 16'h0c68, 16'h0c67, 16'h0c66, 16'h0c65, 16'h0c64},
                                {16'h0c63, 16'h0c62, 16'h0c61, 16'h0c60, 16'h0c5f, 16'h0c5e, 16'h0c5d, 16'h0c5c, 16'h0c5b, 16'h0c5a, 16'h0c59, 16'h0c58, 16'h0c57, 16'h0c56, 16'h0c55, 16'h0c54, 16'h0c53, 16'h0c52, 16'h0c51, 16'h0c50, 16'h0c4f, 16'h0c4e, 16'h0c4d, 16'h0c4c, 16'h0c4b, 16'h0c4a, 16'h0c49, 16'h0c48, 16'h0c47, 16'h0c46, 16'h0c45, 16'h0c44, 16'h0c43, 16'h0c42, 16'h0c41, 16'h0c40, 16'h0c3f, 16'h0c3e, 16'h0c3d, 16'h0c3c, 16'h0c3b, 16'h0c3a, 16'h0c39, 16'h0c38, 16'h0c37, 16'h0c36, 16'h0c35, 16'h0c34, 16'h0c33, 16'h0c32, 16'h0c31, 16'h0c30, 16'h0c2f, 16'h0c2e, 16'h0c2d, 16'h0c2c, 16'h0c2b, 16'h0c2a, 16'h0c29, 16'h0c28, 16'h0c27, 16'h0c26, 16'h0c25, 16'h0c24},
                                {16'h0c23, 16'h0c22, 16'h0c21, 16'h0c20, 16'h0c1f, 16'h0c1e, 16'h0c1d, 16'h0c1c, 16'h0c1b, 16'h0c1a, 16'h0c19, 16'h0c18, 16'h0c17, 16'h0c16, 16'h0c15, 16'h0c14, 16'h0c13, 16'h0c12, 16'h0c11, 16'h0c10, 16'h0c0f, 16'h0c0e, 16'h0c0d, 16'h0c0c, 16'h0c0b, 16'h0c0a, 16'h0c09, 16'h0c08, 16'h0c07, 16'h0c06, 16'h0c05, 16'h0c04, 16'h0c03, 16'h0c02, 16'h0c01, 16'h0c00, 16'h0bff, 16'h0bfe, 16'h0bfd, 16'h0bfc, 16'h0bfb, 16'h0bfa, 16'h0bf9, 16'h0bf8, 16'h0bf7, 16'h0bf6, 16'h0bf5, 16'h0bf4, 16'h0bf3, 16'h0bf2, 16'h0bf1, 16'h0bf0, 16'h0bef, 16'h0bee, 16'h0bed, 16'h0bec, 16'h0beb, 16'h0bea, 16'h0be9, 16'h0be8, 16'h0be7, 16'h0be6, 16'h0be5, 16'h0be4},
                                {16'h0be3, 16'h0be2, 16'h0be1, 16'h0be0, 16'h0bdf, 16'h0bde, 16'h0bdd, 16'h0bdc, 16'h0bdb, 16'h0bda, 16'h0bd9, 16'h0bd8, 16'h0bd7, 16'h0bd6, 16'h0bd5, 16'h0bd4, 16'h0bd3, 16'h0bd2, 16'h0bd1, 16'h0bd0, 16'h0bcf, 16'h0bce, 16'h0bcd, 16'h0bcc, 16'h0bcb, 16'h0bca, 16'h0bc9, 16'h0bc8, 16'h0bc7, 16'h0bc6, 16'h0bc5, 16'h0bc4, 16'h0bc3, 16'h0bc2, 16'h0bc1, 16'h0bc0, 16'h0bbf, 16'h0bbe, 16'h0bbd, 16'h0bbc, 16'h0bbb, 16'h0bba, 16'h0bb9, 16'h0bb8, 16'h0bb7, 16'h0bb6, 16'h0bb5, 16'h0bb4, 16'h0bb3, 16'h0bb2, 16'h0bb1, 16'h0bb0, 16'h0baf, 16'h0bae, 16'h0bad, 16'h0bac, 16'h0bab, 16'h0baa, 16'h0ba9, 16'h0ba8, 16'h0ba7, 16'h0ba6, 16'h0ba5, 16'h0ba4},
                                {16'h0ba3, 16'h0ba2, 16'h0ba1, 16'h0ba0, 16'h0b9f, 16'h0b9e, 16'h0b9d, 16'h0b9c, 16'h0b9b, 16'h0b9a, 16'h0b99, 16'h0b98, 16'h0b97, 16'h0b96, 16'h0b95, 16'h0b94, 16'h0b93, 16'h0b92, 16'h0b91, 16'h0b90, 16'h0b8f, 16'h0b8e, 16'h0b8d, 16'h0b8c, 16'h0b8b, 16'h0b8a, 16'h0b89, 16'h0b88, 16'h0b87, 16'h0b86, 16'h0b85, 16'h0b84, 16'h0b83, 16'h0b82, 16'h0b81, 16'h0b80, 16'h0b7f, 16'h0b7e, 16'h0b7d, 16'h0b7c, 16'h0b7b, 16'h0b7a, 16'h0b79, 16'h0b78, 16'h0b77, 16'h0b76, 16'h0b75, 16'h0b74, 16'h0b73, 16'h0b72, 16'h0b71, 16'h0b70, 16'h0b6f, 16'h0b6e, 16'h0b6d, 16'h0b6c, 16'h0b6b, 16'h0b6a, 16'h0b69, 16'h0b68, 16'h0b67, 16'h0b66, 16'h0b65, 16'h0b64},
                                {16'h0b63, 16'h0b62, 16'h0b61, 16'h0b60, 16'h0b5f, 16'h0b5e, 16'h0b5d, 16'h0b5c, 16'h0b5b, 16'h0b5a, 16'h0b59, 16'h0b58, 16'h0b57, 16'h0b56, 16'h0b55, 16'h0b54, 16'h0b53, 16'h0b52, 16'h0b51, 16'h0b50, 16'h0b4f, 16'h0b4e, 16'h0b4d, 16'h0b4c, 16'h0b4b, 16'h0b4a, 16'h0b49, 16'h0b48, 16'h0b47, 16'h0b46, 16'h0b45, 16'h0b44, 16'h0b43, 16'h0b42, 16'h0b41, 16'h0b40, 16'h0b3f, 16'h0b3e, 16'h0b3d, 16'h0b3c, 16'h0b3b, 16'h0b3a, 16'h0b39, 16'h0b38, 16'h0b37, 16'h0b36, 16'h0b35, 16'h0b34, 16'h0b33, 16'h0b32, 16'h0b31, 16'h0b30, 16'h0b2f, 16'h0b2e, 16'h0b2d, 16'h0b2c, 16'h0b2b, 16'h0b2a, 16'h0b29, 16'h0b28, 16'h0b27, 16'h0b26, 16'h0b25, 16'h0b24},
                                {16'h0b23, 16'h0b22, 16'h0b21, 16'h0b20, 16'h0b1f, 16'h0b1e, 16'h0b1d, 16'h0b1c, 16'h0b1b, 16'h0b1a, 16'h0b19, 16'h0b18, 16'h0b17, 16'h0b16, 16'h0b15, 16'h0b14, 16'h0b13, 16'h0b12, 16'h0b11, 16'h0b10, 16'h0b0f, 16'h0b0e, 16'h0b0d, 16'h0b0c, 16'h0b0b, 16'h0b0a, 16'h0b09, 16'h0b08, 16'h0b07, 16'h0b06, 16'h0b05, 16'h0b04, 16'h0b03, 16'h0b02, 16'h0b01, 16'h0b00, 16'h0aff, 16'h0afe, 16'h0afd, 16'h0afc, 16'h0afb, 16'h0afa, 16'h0af9, 16'h0af8, 16'h0af7, 16'h0af6, 16'h0af5, 16'h0af4, 16'h0af3, 16'h0af2, 16'h0af1, 16'h0af0, 16'h0aef, 16'h0aee, 16'h0aed, 16'h0aec, 16'h0aeb, 16'h0aea, 16'h0ae9, 16'h0ae8, 16'h0ae7, 16'h0ae6, 16'h0ae5, 16'h0ae4},
                                {16'h0ae3, 16'h0ae2, 16'h0ae1, 16'h0ae0, 16'h0adf, 16'h0ade, 16'h0add, 16'h0adc, 16'h0adb, 16'h0ada, 16'h0ad9, 16'h0ad8, 16'h0ad7, 16'h0ad6, 16'h0ad5, 16'h0ad4, 16'h0ad3, 16'h0ad2, 16'h0ad1, 16'h0ad0, 16'h0acf, 16'h0ace, 16'h0acd, 16'h0acc, 16'h0acb, 16'h0aca, 16'h0ac9, 16'h0ac8, 16'h0ac7, 16'h0ac6, 16'h0ac5, 16'h0ac4, 16'h0ac3, 16'h0ac2, 16'h0ac1, 16'h0ac0, 16'h0abf, 16'h0abe, 16'h0abd, 16'h0abc, 16'h0abb, 16'h0aba, 16'h0ab9, 16'h0ab8, 16'h0ab7, 16'h0ab6, 16'h0ab5, 16'h0ab4, 16'h0ab3, 16'h0ab2, 16'h0ab1, 16'h0ab0, 16'h0aaf, 16'h0aae, 16'h0aad, 16'h0aac, 16'h0aab, 16'h0aaa, 16'h0aa9, 16'h0aa8, 16'h0aa7, 16'h0aa6, 16'h0aa5, 16'h0aa4},
                                {16'h0aa3, 16'h0aa2, 16'h0aa1, 16'h0aa0, 16'h0a9f, 16'h0a9e, 16'h0a9d, 16'h0a9c, 16'h0a9b, 16'h0a9a, 16'h0a99, 16'h0a98, 16'h0a97, 16'h0a96, 16'h0a95, 16'h0a94, 16'h0a93, 16'h0a92, 16'h0a91, 16'h0a90, 16'h0a8f, 16'h0a8e, 16'h0a8d, 16'h0a8c, 16'h0a8b, 16'h0a8a, 16'h0a89, 16'h0a88, 16'h0a87, 16'h0a86, 16'h0a85, 16'h0a84, 16'h0a83, 16'h0a82, 16'h0a81, 16'h0a80, 16'h0a7f, 16'h0a7e, 16'h0a7d, 16'h0a7c, 16'h0a7b, 16'h0a7a, 16'h0a79, 16'h0a78, 16'h0a77, 16'h0a76, 16'h0a75, 16'h0a74, 16'h0a73, 16'h0a72, 16'h0a71, 16'h0a70, 16'h0a6f, 16'h0a6e, 16'h0a6d, 16'h0a6c, 16'h0a6b, 16'h0a6a, 16'h0a69, 16'h0a68, 16'h0a67, 16'h0a66, 16'h0a65, 16'h0a64},
                                {16'h0a63, 16'h0a62, 16'h0a61, 16'h0a60, 16'h0a5f, 16'h0a5e, 16'h0a5d, 16'h0a5c, 16'h0a5b, 16'h0a5a, 16'h0a59, 16'h0a58, 16'h0a57, 16'h0a56, 16'h0a55, 16'h0a54, 16'h0a53, 16'h0a52, 16'h0a51, 16'h0a50, 16'h0a4f, 16'h0a4e, 16'h0a4d, 16'h0a4c, 16'h0a4b, 16'h0a4a, 16'h0a49, 16'h0a48, 16'h0a47, 16'h0a46, 16'h0a45, 16'h0a44, 16'h0a43, 16'h0a42, 16'h0a41, 16'h0a40, 16'h0a3f, 16'h0a3e, 16'h0a3d, 16'h0a3c, 16'h0a3b, 16'h0a3a, 16'h0a39, 16'h0a38, 16'h0a37, 16'h0a36, 16'h0a35, 16'h0a34, 16'h0a33, 16'h0a32, 16'h0a31, 16'h0a30, 16'h0a2f, 16'h0a2e, 16'h0a2d, 16'h0a2c, 16'h0a2b, 16'h0a2a, 16'h0a29, 16'h0a28, 16'h0a27, 16'h0a26, 16'h0a25, 16'h0a24},
                                {16'h0a23, 16'h0a22, 16'h0a21, 16'h0a20, 16'h0a1f, 16'h0a1e, 16'h0a1d, 16'h0a1c, 16'h0a1b, 16'h0a1a, 16'h0a19, 16'h0a18, 16'h0a17, 16'h0a16, 16'h0a15, 16'h0a14, 16'h0a13, 16'h0a12, 16'h0a11, 16'h0a10, 16'h0a0f, 16'h0a0e, 16'h0a0d, 16'h0a0c, 16'h0a0b, 16'h0a0a, 16'h0a09, 16'h0a08, 16'h0a07, 16'h0a06, 16'h0a05, 16'h0a04, 16'h0a03, 16'h0a02, 16'h0a01, 16'h0a00, 16'h09ff, 16'h09fe, 16'h09fd, 16'h09fc, 16'h09fb, 16'h09fa, 16'h09f9, 16'h09f8, 16'h09f7, 16'h09f6, 16'h09f5, 16'h09f4, 16'h09f3, 16'h09f2, 16'h09f1, 16'h09f0, 16'h09ef, 16'h09ee, 16'h09ed, 16'h09ec, 16'h09eb, 16'h09ea, 16'h09e9, 16'h09e8, 16'h09e7, 16'h09e6, 16'h09e5, 16'h09e4},
                                {16'h09e3, 16'h09e2, 16'h09e1, 16'h09e0, 16'h09df, 16'h09de, 16'h09dd, 16'h09dc, 16'h09db, 16'h09da, 16'h09d9, 16'h09d8, 16'h09d7, 16'h09d6, 16'h09d5, 16'h09d4, 16'h09d3, 16'h09d2, 16'h09d1, 16'h09d0, 16'h09cf, 16'h09ce, 16'h09cd, 16'h09cc, 16'h09cb, 16'h09ca, 16'h09c9, 16'h09c8, 16'h09c7, 16'h09c6, 16'h09c5, 16'h09c4, 16'h09c3, 16'h09c2, 16'h09c1, 16'h09c0, 16'h09bf, 16'h09be, 16'h09bd, 16'h09bc, 16'h09bb, 16'h09ba, 16'h09b9, 16'h09b8, 16'h09b7, 16'h09b6, 16'h09b5, 16'h09b4, 16'h09b3, 16'h09b2, 16'h09b1, 16'h09b0, 16'h09af, 16'h09ae, 16'h09ad, 16'h09ac, 16'h09ab, 16'h09aa, 16'h09a9, 16'h09a8, 16'h09a7, 16'h09a6, 16'h09a5, 16'h09a4},
                                {16'h09a3, 16'h09a2, 16'h09a1, 16'h09a0, 16'h099f, 16'h099e, 16'h099d, 16'h099c, 16'h099b, 16'h099a, 16'h0999, 16'h0998, 16'h0997, 16'h0996, 16'h0995, 16'h0994, 16'h0993, 16'h0992, 16'h0991, 16'h0990, 16'h098f, 16'h098e, 16'h098d, 16'h098c, 16'h098b, 16'h098a, 16'h0989, 16'h0988, 16'h0987, 16'h0986, 16'h0985, 16'h0984, 16'h0983, 16'h0982, 16'h0981, 16'h0980, 16'h097f, 16'h097e, 16'h097d, 16'h097c, 16'h097b, 16'h097a, 16'h0979, 16'h0978, 16'h0977, 16'h0976, 16'h0975, 16'h0974, 16'h0973, 16'h0972, 16'h0971, 16'h0970, 16'h096f, 16'h096e, 16'h096d, 16'h096c, 16'h096b, 16'h096a, 16'h0969, 16'h0968, 16'h0967, 16'h0966, 16'h0965, 16'h0964},
                                {16'h0963, 16'h0962, 16'h0961, 16'h0960, 16'h095f, 16'h095e, 16'h095d, 16'h095c, 16'h095b, 16'h095a, 16'h0959, 16'h0958, 16'h0957, 16'h0956, 16'h0955, 16'h0954, 16'h0953, 16'h0952, 16'h0951, 16'h0950, 16'h094f, 16'h094e, 16'h094d, 16'h094c, 16'h094b, 16'h094a, 16'h0949, 16'h0948, 16'h0947, 16'h0946, 16'h0945, 16'h0944, 16'h0943, 16'h0942, 16'h0941, 16'h0940, 16'h093f, 16'h093e, 16'h093d, 16'h093c, 16'h093b, 16'h093a, 16'h0939, 16'h0938, 16'h0937, 16'h0936, 16'h0935, 16'h0934, 16'h0933, 16'h0932, 16'h0931, 16'h0930, 16'h092f, 16'h092e, 16'h092d, 16'h092c, 16'h092b, 16'h092a, 16'h0929, 16'h0928, 16'h0927, 16'h0926, 16'h0925, 16'h0924},
                                {16'h0923, 16'h0922, 16'h0921, 16'h0920, 16'h091f, 16'h091e, 16'h091d, 16'h091c, 16'h091b, 16'h091a, 16'h0919, 16'h0918, 16'h0917, 16'h0916, 16'h0915, 16'h0914, 16'h0913, 16'h0912, 16'h0911, 16'h0910, 16'h090f, 16'h090e, 16'h090d, 16'h090c, 16'h090b, 16'h090a, 16'h0909, 16'h0908, 16'h0907, 16'h0906, 16'h0905, 16'h0904, 16'h0903, 16'h0902, 16'h0901, 16'h0900, 16'h08ff, 16'h08fe, 16'h08fd, 16'h08fc, 16'h08fb, 16'h08fa, 16'h08f9, 16'h08f8, 16'h08f7, 16'h08f6, 16'h08f5, 16'h08f4, 16'h08f3, 16'h08f2, 16'h08f1, 16'h08f0, 16'h08ef, 16'h08ee, 16'h08ed, 16'h08ec, 16'h08eb, 16'h08ea, 16'h08e9, 16'h08e8, 16'h08e7, 16'h08e6, 16'h08e5, 16'h08e4},
                                {16'h08e3, 16'h08e2, 16'h08e1, 16'h08e0, 16'h08df, 16'h08de, 16'h08dd, 16'h08dc, 16'h08db, 16'h08da, 16'h08d9, 16'h08d8, 16'h08d7, 16'h08d6, 16'h08d5, 16'h08d4, 16'h08d3, 16'h08d2, 16'h08d1, 16'h08d0, 16'h08cf, 16'h08ce, 16'h08cd, 16'h08cc, 16'h08cb, 16'h08ca, 16'h08c9, 16'h08c8, 16'h08c7, 16'h08c6, 16'h08c5, 16'h08c4, 16'h08c3, 16'h08c2, 16'h08c1, 16'h08c0, 16'h08bf, 16'h08be, 16'h08bd, 16'h08bc, 16'h08bb, 16'h08ba, 16'h08b9, 16'h08b8, 16'h08b7, 16'h08b6, 16'h08b5, 16'h08b4, 16'h08b3, 16'h08b2, 16'h08b1, 16'h08b0, 16'h08af, 16'h08ae, 16'h08ad, 16'h08ac, 16'h08ab, 16'h08aa, 16'h08a9, 16'h08a8, 16'h08a7, 16'h08a6, 16'h08a5, 16'h08a4},
                                {16'h08a3, 16'h08a2, 16'h08a1, 16'h08a0, 16'h089f, 16'h089e, 16'h089d, 16'h089c, 16'h089b, 16'h089a, 16'h089a, 16'h089a, 16'h089a, 16'h089a, 16'h08a1, 16'h08aa, 16'h08b3, 16'h08bc, 16'h08c5, 16'h08ce, 16'h08d7, 16'h08e0, 16'h08e9, 16'h08f2, 16'h08fb, 16'h0904, 16'h090d, 16'h0916, 16'h091f, 16'h0928, 16'h0931, 16'h093a, 16'h0943, 16'h094c, 16'h0955, 16'h095e, 16'h0967, 16'h0970, 16'h0979, 16'h0982, 16'h098b, 16'h0994, 16'h099d, 16'h09a6, 16'h09af, 16'h09b8, 16'h09c1, 16'h09ca, 16'h09d3, 16'h09dc, 16'h09e5, 16'h09ee, 16'h09f7, 16'h0a00, 16'h0a09, 16'h0a12, 16'h0a1b, 16'h0a24, 16'h0a2d, 16'h0a36, 16'h0a3f, 16'h0a48, 16'h0a51, 16'h0a5a},
                                {16'h0a63, 16'h0a6c, 16'h0a75, 16'h0a7e, 16'h0a87, 16'h0a90, 16'h0a99, 16'h0aa2, 16'h0aab, 16'h0ab4, 16'h0abd, 16'h0ac6, 16'h0acf, 16'h0ad8, 16'h0ae1, 16'h0aea, 16'h0af3, 16'h0afc, 16'h0b05, 16'h0b0e, 16'h0b17, 16'h0b20, 16'h0b29, 16'h0b32, 16'h0b3b, 16'h0b44, 16'h0b4d, 16'h0b56, 16'h0b5f, 16'h0b68, 16'h0b71, 16'h0b7a, 16'h0b83, 16'h0b8c, 16'h0b95, 16'h0b9e, 16'h0ba7, 16'h0bb0, 16'h0bb9, 16'h0bc2, 16'h0bcb, 16'h0bd4, 16'h0bdd, 16'h0be6, 16'h0bef, 16'h0bf8, 16'h0c01, 16'h0c0a, 16'h0c13, 16'h0c1c, 16'h0c25, 16'h0c2e, 16'h0c37, 16'h0c40, 16'h0c49, 16'h0c52, 16'h0c5b, 16'h0c64, 16'h0c6d, 16'h0c76, 16'h0c7f, 16'h0c88, 16'h0c91, 16'h0c9a},
                                {16'h0ca3, 16'h0cac, 16'h0cb5, 16'h0cbe, 16'h0cc7, 16'h0cd0, 16'h0cd9, 16'h0ce2, 16'h0ceb, 16'h0cf4, 16'h0cfd, 16'h0d06, 16'h0d0f, 16'h0d18, 16'h0d21, 16'h0d2a, 16'h0d33, 16'h0d3c, 16'h0d45, 16'h0d4e, 16'h0d57, 16'h0d60, 16'h0d69, 16'h0d72, 16'h0d7b, 16'h0d84, 16'h0d8d, 16'h0d96, 16'h0d9f, 16'h0da8, 16'h0db1, 16'h0dba, 16'h0dc3, 16'h0dcc, 16'h0dd5, 16'h0dde, 16'h0de7, 16'h0df0, 16'h0df9, 16'h0e02, 16'h0e0b, 16'h0e14, 16'h0e1d, 16'h0e26, 16'h0e2f, 16'h0e38, 16'h0e41, 16'h0e4a, 16'h0e53, 16'h0e5c, 16'h0e65, 16'h0e6e, 16'h0e77, 16'h0e80, 16'h0e89, 16'h0e92, 16'h0e9b, 16'h0ea4, 16'h0ead, 16'h0eb6, 16'h0ebf, 16'h0ec8, 16'h0ed1, 16'h0eda},
                                {16'h0ee3, 16'h0eec, 16'h0ef5, 16'h0efe, 16'h0f07, 16'h0f10, 16'h0f19, 16'h0f22, 16'h0f2b, 16'h0f34, 16'h0f3d, 16'h0f46, 16'h0f4f, 16'h0f58, 16'h0f61, 16'h0f6a, 16'h0f73, 16'h0f7c, 16'h0f85, 16'h0f8e, 16'h0f97, 16'h0fa0, 16'h0fa9, 16'h0fb2, 16'h0fbb, 16'h0fc4, 16'h0fcd, 16'h0fd6, 16'h0fdf, 16'h0fe8, 16'h0ff1, 16'h0ffa, 16'h1003, 16'h100c, 16'h1015, 16'h101e, 16'h1027, 16'h1030, 16'h1039, 16'h1042, 16'h104b, 16'h1054, 16'h105d, 16'h1071, 16'h1079, 16'h1081, 16'h1089, 16'h1091, 16'h1099, 16'h10a1, 16'h10a9, 16'h10b1, 16'h10b9, 16'h10c1, 16'h10c9, 16'h10d1, 16'h10d9, 16'h10e1, 16'h10e9, 16'h10f1, 16'h10f9, 16'h1101, 16'h1109, 16'h1111},
                                {16'h1119, 16'h1121, 16'h1129, 16'h1131, 16'h1139, 16'h1141, 16'h1149, 16'h1151, 16'h1159, 16'h1161, 16'h1169, 16'h1171, 16'h1179, 16'h1181, 16'h1189, 16'h1191, 16'h1199, 16'h11a1, 16'h11a9, 16'h11b1, 16'h11b9, 16'h11c1, 16'h11c9, 16'h11d1, 16'h11d9, 16'h11e1, 16'h11e9, 16'h11f1, 16'h11f9, 16'h1201, 16'h1209, 16'h1211, 16'h1219, 16'h1221, 16'h1229, 16'h1231, 16'h1239, 16'h1241, 16'h1249, 16'h1251, 16'h1259, 16'h1261, 16'h1269, 16'h1271, 16'h1279, 16'h1281, 16'h1289, 16'h1291, 16'h1299, 16'h12a1, 16'h12a9, 16'h12b1, 16'h12b9, 16'h12c1, 16'h12c9, 16'h12d1, 16'h12d9, 16'h12e1, 16'h12e9, 16'h12f1, 16'h12f9, 16'h1301, 16'h1309, 16'h1311},
                                {16'h1319, 16'h1321, 16'h1329, 16'h1331, 16'h1339, 16'h1341, 16'h1349, 16'h1351, 16'h1359, 16'h1361, 16'h1369, 16'h1371, 16'h1379, 16'h1381, 16'h1389, 16'h1391, 16'h1399, 16'h13a1, 16'h13a9, 16'h13b1, 16'h13b9, 16'h13c1, 16'h13c9, 16'h13d1, 16'h13d9, 16'h13e1, 16'h13e9, 16'h13f1, 16'h13f9, 16'h1401, 16'h1409, 16'h1411, 16'h1419, 16'h1421, 16'h1429, 16'h1431, 16'h1439, 16'h1441, 16'h1449, 16'h1451, 16'h1459, 16'h1461, 16'h1469, 16'h1471, 16'h1479, 16'h1481, 16'h1489, 16'h1491, 16'h1499, 16'h14a1, 16'h14a9, 16'h14b1, 16'h14b9, 16'h14c1, 16'h14c9, 16'h14d1, 16'h14d9, 16'h14e1, 16'h14e9, 16'h14f1, 16'h14f9, 16'h1501, 16'h1509, 16'h1511},
                                {16'h1519, 16'h1521, 16'h1529, 16'h1531, 16'h1539, 16'h1541, 16'h1549, 16'h1551, 16'h1559, 16'h1561, 16'h1569, 16'h1571, 16'h1579, 16'h1581, 16'h1589, 16'h1591, 16'h1599, 16'h15a1, 16'h15a9, 16'h15b1, 16'h15b9, 16'h15c1, 16'h15c9, 16'h15d1, 16'h15d9, 16'h15e1, 16'h15e9, 16'h15f1, 16'h15f9, 16'h1601, 16'h1609, 16'h1611, 16'h1619, 16'h1621, 16'h1629, 16'h1631, 16'h1639, 16'h1641, 16'h1649, 16'h1651, 16'h1659, 16'h1661, 16'h1669, 16'h1671, 16'h1679, 16'h1681, 16'h1689, 16'h1691, 16'h1699, 16'h16a1, 16'h16a9, 16'h16b1, 16'h16b9, 16'h16c1, 16'h16c9, 16'h16d1, 16'h16d9, 16'h16e1, 16'h16e9, 16'h16f1, 16'h16f9, 16'h1701, 16'h1709, 16'h1711},
                                {16'h1719, 16'h1721, 16'h1729, 16'h1731, 16'h1739, 16'h1741, 16'h1749, 16'h1751, 16'h1759, 16'h1761, 16'h1769, 16'h1771, 16'h1779, 16'h1781, 16'h1789, 16'h1791, 16'h1799, 16'h17a1, 16'h17a9, 16'h17b1, 16'h17b9, 16'h17c1, 16'h17c9, 16'h17d1, 16'h17d9, 16'h17e1, 16'h17e9, 16'h17f1, 16'h17f9, 16'h1801, 16'h1809, 16'h1811, 16'h1819, 16'h1821, 16'h1829, 16'h1831, 16'h1839, 16'h1841, 16'h1849, 16'h1851, 16'h1859, 16'h1861, 16'h1869, 16'h1871, 16'h1879, 16'h1881, 16'h1889, 16'h1891, 16'h1899, 16'h18a1, 16'h18a9, 16'h18ad, 16'h18be, 16'h18cf, 16'h18e0, 16'h18f1, 16'h1902, 16'h1913, 16'h1924, 16'h1935, 16'h1946, 16'h1957, 16'h1968, 16'h1979},
                                {16'h198a, 16'h199b, 16'h19ac, 16'h19bd, 16'h19ce, 16'h19df, 16'h19f0, 16'h1a01, 16'h1a12, 16'h1a23, 16'h1a34, 16'h1a45, 16'h1a56, 16'h1a67, 16'h1a78, 16'h1a89, 16'h1a9a, 16'h1aab, 16'h1abc, 16'h1acd, 16'h1ade, 16'h1aef, 16'h1b00, 16'h1b11, 16'h1b22, 16'h1b33, 16'h1b44, 16'h1b55, 16'h1b66, 16'h1b77, 16'h1b88, 16'h1b99, 16'h1baa, 16'h1bbb, 16'h1bcc, 16'h1bdd, 16'h1bee, 16'h1bff, 16'h1c10, 16'h1c21, 16'h1c32, 16'h1c43, 16'h1c54, 16'h1c65, 16'h1c76, 16'h1c87, 16'h1c98, 16'h1ca9, 16'h1cba, 16'h1ccb, 16'h1cdc, 16'h1ced, 16'h1cfe, 16'h1d0f, 16'h1d20, 16'h1d31, 16'h1d42, 16'h1d53, 16'h1d64, 16'h1d75, 16'h1d86, 16'h1d97, 16'h1da8, 16'h1db9},
                                {16'h1dca, 16'h1ddb, 16'h1dec, 16'h1dfd, 16'h1e0e, 16'h1e1f, 16'h1e30, 16'h1e41, 16'h1e52, 16'h1e63, 16'h1e74, 16'h1e85, 16'h1e96, 16'h1ea7, 16'h1eb8, 16'h1ec9, 16'h1eda, 16'h1eeb, 16'h1efc, 16'h1f0d, 16'h1f1e, 16'h1f2f, 16'h1f40, 16'h1f51, 16'h1f62, 16'h1f73, 16'h1f84, 16'h1f95, 16'h1fa6, 16'h1fb7, 16'h1fc8, 16'h1fd9, 16'h1fea, 16'h1ffb, 16'h200c, 16'h201d, 16'h201d, 16'h201d, 16'h201d, 16'h201f, 16'h202e, 16'h203d, 16'h204c, 16'h205b, 16'h206a, 16'h2079, 16'h2088, 16'h2097, 16'h20a6, 16'h20b5, 16'h20c4, 16'h20d3, 16'h20e2, 16'h20f1, 16'h2100, 16'h210f, 16'h211e, 16'h212d, 16'h213c, 16'h214b, 16'h215a, 16'h2169, 16'h2178, 16'h2187},
                                {16'h2196, 16'h21a5, 16'h21b4, 16'h21c3, 16'h21d2, 16'h21e1, 16'h21f0, 16'h21ff, 16'h220e, 16'h221d, 16'h222c, 16'h223b, 16'h224a, 16'h2259, 16'h2268, 16'h2277, 16'h2286, 16'h2295, 16'h22a4, 16'h22b3, 16'h22c2, 16'h22d1, 16'h22e0, 16'h22ef, 16'h22fe, 16'h230d, 16'h231c, 16'h232b, 16'h233a, 16'h2349, 16'h2358, 16'h2367, 16'h2376, 16'h2385, 16'h2394, 16'h23a3, 16'h23b2, 16'h23c1, 16'h23d0, 16'h23df, 16'h23ee, 16'h23fd, 16'h240c, 16'h241b, 16'h242a, 16'h2439, 16'h2448, 16'h2457, 16'h2466, 16'h2475, 16'h2484, 16'h2493, 16'h24a2, 16'h24b1, 16'h24c0, 16'h24cf, 16'h24de, 16'h24ed, 16'h24fc, 16'h250b, 16'h251a, 16'h2529, 16'h2538, 16'h2547},
                                {16'h2556, 16'h2565, 16'h2574, 16'h2583, 16'h2592, 16'h25a1, 16'h25b0, 16'h25bf, 16'h25ce, 16'h25dd, 16'h25ec, 16'h25fb, 16'h260a, 16'h2619, 16'h2628, 16'h2637, 16'h2646, 16'h2655, 16'h2664, 16'h2673, 16'h2682, 16'h2691, 16'h26a0, 16'h26af, 16'h26be, 16'h26cd, 16'h26dc, 16'h26eb, 16'h26fa, 16'h2709, 16'h2718, 16'h2727, 16'h2736, 16'h2745, 16'h2754, 16'h2763, 16'h2772, 16'h2781, 16'h2790, 16'h299b, 16'h299c, 16'h299d, 16'h299e, 16'h299f, 16'h29a0, 16'h29a1, 16'h29a2, 16'h29a3, 16'h29a4, 16'h29a5, 16'h29a6, 16'h29a7, 16'h29a8, 16'h29a9, 16'h29aa, 16'h29ab, 16'h29ac, 16'h29ad, 16'h29ae, 16'h29af, 16'h29b0, 16'h29b1, 16'h29b2, 16'h29b3},
                                {16'h29b4, 16'h29b5, 16'h29b6, 16'h29b7, 16'h29b8, 16'h29b9, 16'h29ba, 16'h29bb, 16'h29bc, 16'h29bd, 16'h29be, 16'h29bf, 16'h29c0, 16'h29c1, 16'h29c2, 16'h29c3, 16'h29c4, 16'h29c5, 16'h29c6, 16'h29c7, 16'h29c8, 16'h29c9, 16'h29ca, 16'h29cb, 16'h29cc, 16'h29cd, 16'h29ce, 16'h29cf, 16'h29d0, 16'h29d1, 16'h29d2, 16'h29d3, 16'h29d4, 16'h29d5, 16'h29d6, 16'h29d7, 16'h29d8, 16'h29d9, 16'h29da, 16'h29db, 16'h29dc, 16'h29dd, 16'h29de, 16'h29df, 16'h29e0, 16'h29e1, 16'h29e2, 16'h29e3, 16'h29e4, 16'h29e5, 16'h29e6, 16'h29e7, 16'h29e8, 16'h29e9, 16'h29ea, 16'h29eb, 16'h29ec, 16'h29ed, 16'h29ee, 16'h29ef, 16'h29f0, 16'h29f1, 16'h29f2, 16'h29f3},
                                {16'h29f4, 16'h29f5, 16'h29f6, 16'h29f7, 16'h29f8, 16'h29f9, 16'h29fa, 16'h29fb, 16'h29fc, 16'h29fd, 16'h29fe, 16'h29ff, 16'h2a00, 16'h2a01, 16'h2a02, 16'h2a03, 16'h2a04, 16'h2a05, 16'h2a06, 16'h2a07, 16'h2a08, 16'h2a09, 16'h2a0a, 16'h2a0b, 16'h2a0c, 16'h2a0d, 16'h2a0e, 16'h2a0f, 16'h2a10, 16'h2a11, 16'h2a12, 16'h2a13, 16'h2a14, 16'h2a15, 16'h2a16, 16'h2a17, 16'h2a18, 16'h2a19, 16'h2a1a, 16'h2a1b, 16'h2a1c, 16'h2a1d, 16'h2a1e, 16'h2a1f, 16'h2a20, 16'h2a21, 16'h2a22, 16'h2a23, 16'h2a24, 16'h2a25, 16'h2a26, 16'h2a27, 16'h2a28, 16'h2a29, 16'h2a2a, 16'h2a2b, 16'h2a2c, 16'h2a2d, 16'h2a2e, 16'h2a2f, 16'h2a30, 16'h2a31, 16'h2a32, 16'h2a33},
                                {16'h2a34, 16'h2a35, 16'h2a36, 16'h2a37, 16'h2a38, 16'h2a39, 16'h2a3a, 16'h2a3b, 16'h2a3c, 16'h2a3d, 16'h2a3e, 16'h2a3f, 16'h2a40, 16'h2a41, 16'h2a42, 16'h2a43, 16'h2a44, 16'h2a45, 16'h2a46, 16'h2a47, 16'h2a48, 16'h2a49, 16'h2a4a, 16'h2a4b, 16'h2a4c, 16'h2a4d, 16'h2a4e, 16'h2a4f, 16'h2a50, 16'h2a51, 16'h2a52, 16'h2a53, 16'h2a54, 16'h2a55, 16'h2a56, 16'h2a57, 16'h2a58, 16'h2a59, 16'h2a5a, 16'h2a5b, 16'h2a5c, 16'h2a5d, 16'h2a5e, 16'h2a5f, 16'h2a60, 16'h2a61, 16'h2a62, 16'h2a63, 16'h2a64, 16'h2a65, 16'h2a66, 16'h2a67, 16'h2a68, 16'h2a69, 16'h2a6a, 16'h2a6b, 16'h2a6c, 16'h2a6d, 16'h2a6e, 16'h2a6f, 16'h2a70, 16'h2a71, 16'h2a72, 16'h2a73},
                                {16'h2a74, 16'h2a75, 16'h2a76, 16'h2a77, 16'h2a78, 16'h2a79, 16'h2a7a, 16'h2a7b, 16'h2a7c, 16'h2a7d, 16'h2a7e, 16'h2a7f, 16'h2a80, 16'h2a81, 16'h2a82, 16'h2a83, 16'h2a84, 16'h2a85, 16'h2a86, 16'h2a87, 16'h2a88, 16'h2a89, 16'h2a8a, 16'h2a8b, 16'h2a8c, 16'h2a8d, 16'h2a8e, 16'h2a8f, 16'h2a90, 16'h2a91, 16'h2a92, 16'h2a93, 16'h2a94, 16'h2a95, 16'h2a96, 16'h2a97, 16'h2a98, 16'h2a99, 16'h2a9a, 16'h2a9b, 16'h2a9c, 16'h2a9d, 16'h2a9e, 16'h2a9f, 16'h2aa0, 16'h2aa1, 16'h2aa2, 16'h2aa3, 16'h2aa4, 16'h2aa5, 16'h2aa6, 16'h2aa7, 16'h2aa8, 16'h2aa9, 16'h2aaa, 16'h2aab, 16'h2aac, 16'h2aad, 16'h2aae, 16'h2aaf, 16'h2ab0, 16'h2ab1, 16'h2ab2, 16'h2ab3},
                                {16'h2ab4, 16'h2ab5, 16'h2ab6, 16'h2ab7, 16'h2ab8, 16'h2ab9, 16'h2aba, 16'h2abb, 16'h2abc, 16'h2abd, 16'h2abe, 16'h2abf, 16'h2ac0, 16'h2ac1, 16'h2ac2, 16'h2ac3, 16'h2ac4, 16'h2ac5, 16'h2ac6, 16'h2ac7, 16'h2ac8, 16'h2ac9, 16'h2aca, 16'h2acb, 16'h2acc, 16'h2acd, 16'h2ace, 16'h2acf, 16'h2ad0, 16'h2ad1, 16'h2ad2, 16'h2ad3, 16'h2ad4, 16'h2ad5, 16'h2ad6, 16'h2ad7, 16'h2ad8, 16'h2ad9, 16'h2ada, 16'h2adb, 16'h2adc, 16'h2add, 16'h2ade, 16'h2adf, 16'h2ae0, 16'h2ae1, 16'h2ae2, 16'h2ae3, 16'h2ae4, 16'h2ae5, 16'h2ae6, 16'h2ae7, 16'h2ae8, 16'h2ae9, 16'h2aea, 16'h2aeb, 16'h2aec, 16'h2aed, 16'h2aee, 16'h2aef, 16'h2af0, 16'h2af1, 16'h2af2, 16'h2af3},
                                {16'h2af4, 16'h2af5, 16'h2af6, 16'h2af7, 16'h2af8, 16'h2af9, 16'h2afa, 16'h2afb, 16'h2afc, 16'h2afd, 16'h2afe, 16'h2aff, 16'h2b00, 16'h2b01, 16'h2b02, 16'h2b03, 16'h2b04, 16'h2b05, 16'h2b06, 16'h2b07, 16'h2b08, 16'h2b09, 16'h2b0a, 16'h2b0b, 16'h2b0c, 16'h2b0d, 16'h2b0e, 16'h2b0f, 16'h2b10, 16'h2b11, 16'h2b12, 16'h2b13, 16'h2b14, 16'h2b15, 16'h2b16, 16'h2b17, 16'h2b18, 16'h2b19, 16'h2b1a, 16'h2b1b, 16'h2b1c, 16'h2b1d, 16'h2b1e, 16'h2b1f, 16'h2b20, 16'h2b21, 16'h2b22, 16'h2b23, 16'h2b24, 16'h2b25, 16'h2b26, 16'h2b27, 16'h2b28, 16'h2b29, 16'h2b2a, 16'h2b2b, 16'h2b2c, 16'h2b2d, 16'h2b2e, 16'h2b2f, 16'h2b30, 16'h2b31, 16'h2b32, 16'h2b33},
                                {16'h2b34, 16'h2b35, 16'h2b36, 16'h2b37, 16'h2b38, 16'h2b39, 16'h2b3a, 16'h2b3b, 16'h2b3c, 16'h2b3d, 16'h2b3e, 16'h2b3f, 16'h2b40, 16'h2b41, 16'h2b42, 16'h2b43, 16'h2b44, 16'h2b45, 16'h2b46, 16'h2b47, 16'h2b48, 16'h2b49, 16'h2b4a, 16'h2b4b, 16'h2b4c, 16'h2b4d, 16'h2b4e, 16'h2b4f, 16'h2b50, 16'h2b51, 16'h2b52, 16'h2b53, 16'h2b54, 16'h2b55, 16'h2b56, 16'h2b57, 16'h2b58, 16'h2b59, 16'h2b5a, 16'h2b5b, 16'h2b5c, 16'h2b5d, 16'h2b5e, 16'h2b5f, 16'h2b60, 16'h2b61, 16'h2b62, 16'h2b63, 16'h2b64, 16'h2b65, 16'h2b66, 16'h2b67, 16'h2b68, 16'h2b69, 16'h2b6a, 16'h2b6b, 16'h2b6c, 16'h2b6d, 16'h2b6e, 16'h2b6f, 16'h2b70, 16'h2b71, 16'h2b72, 16'h2b73},
                                {16'h2b74, 16'h2b75, 16'h2b76, 16'h2b77, 16'h2b78, 16'h2b79, 16'h2b7a, 16'h2b7b, 16'h2b7c, 16'h2b7d, 16'h2b7e, 16'h2b7f, 16'h2b80, 16'h2b81, 16'h2b82, 16'h2b83, 16'h2b84, 16'h2b85, 16'h2b86, 16'h2b87, 16'h2b88, 16'h2b89, 16'h2b8a, 16'h2b8b, 16'h2b8c, 16'h2b8d, 16'h2b8e, 16'h2b8f, 16'h2b90, 16'h2b91, 16'h2b92, 16'h2b93, 16'h2b94, 16'h2b95, 16'h2b96, 16'h2b97, 16'h2b98, 16'h2b99, 16'h2b9a, 16'h2b9b, 16'h2b9c, 16'h2b9d, 16'h2b9e, 16'h2b9f, 16'h2ba0, 16'h2ba1, 16'h2ba2, 16'h2ba3, 16'h2ba4, 16'h2ba5, 16'h2ba6, 16'h2ba7, 16'h2ba8, 16'h2ba9, 16'h2baa, 16'h2bab, 16'h2bac, 16'h2bad, 16'h2bae, 16'h2baf, 16'h2bb0, 16'h2bb1, 16'h2bb2, 16'h2bb3},
                                {16'h2bb4, 16'h2bb5, 16'h2bb6, 16'h2bb7, 16'h2bb8, 16'h2bb9, 16'h2bba, 16'h2bbb, 16'h2bbc, 16'h2bbd, 16'h2bbe, 16'h2bbf, 16'h2bc0, 16'h2bc1, 16'h2bc2, 16'h2bc3, 16'h2bc4, 16'h2bc5, 16'h2bc6, 16'h2bc7, 16'h2bc8, 16'h2bc9, 16'h2bca, 16'h2bcb, 16'h2bcc, 16'h2bcd, 16'h2bce, 16'h2bcf, 16'h2bd0, 16'h2bd1, 16'h2bd2, 16'h2bd3, 16'h2bd4, 16'h2bd5, 16'h2bd6, 16'h2bd7, 16'h2bd8, 16'h2bd9, 16'h2bda, 16'h2bdb, 16'h2bdc, 16'h2bdd, 16'h2bde, 16'h2bdf, 16'h2be0, 16'h2be1, 16'h2be2, 16'h2be3, 16'h2be4, 16'h2be5, 16'h2be6, 16'h2be7, 16'h2be8, 16'h2be9, 16'h2bea, 16'h2beb, 16'h2bec, 16'h2bed, 16'h2bee, 16'h2bef, 16'h2bf0, 16'h2bf1, 16'h2bf2, 16'h2bf3},
                                {16'h2bf4, 16'h2bf5, 16'h2bf6, 16'h2bf7, 16'h2bf8, 16'h2bf9, 16'h2bfa, 16'h2bfb, 16'h2bfc, 16'h2bfd, 16'h2bfe, 16'h2bff, 16'h2c00, 16'h2c01, 16'h2c02, 16'h2c03, 16'h2c04, 16'h2c05, 16'h2c06, 16'h2c07, 16'h2c08, 16'h2c09, 16'h2c0a, 16'h2c0b, 16'h2c0c, 16'h2c0d, 16'h2c0e, 16'h2c0f, 16'h2c10, 16'h2c11, 16'h2c12, 16'h2c13, 16'h2c14, 16'h2c15, 16'h2c16, 16'h2c17, 16'h2c18, 16'h2c19, 16'h2c1a, 16'h2c1b, 16'h2c1c, 16'h2c1d, 16'h2c1e, 16'h2c1f, 16'h2c20, 16'h2c21, 16'h2c22, 16'h2c23, 16'h2c24, 16'h2c25, 16'h2c26, 16'h2c27, 16'h2c28, 16'h2c29, 16'h2c2a, 16'h2c2b, 16'h2c2c, 16'h2c2d, 16'h2c2e, 16'h2c2f, 16'h2c30, 16'h2c31, 16'h2c32, 16'h2c33},
                                {16'h2c34, 16'h2c35, 16'h2c36, 16'h2c37, 16'h2c38, 16'h2c39, 16'h2c3a, 16'h2c3b, 16'h2c3c, 16'h2c3d, 16'h2c3e, 16'h2c3f, 16'h2c40, 16'h2c41, 16'h2c42, 16'h2c43, 16'h2c44, 16'h2c45, 16'h2c46, 16'h2c47, 16'h2c48, 16'h2c49, 16'h2c4a, 16'h2c4b, 16'h2c4c, 16'h2c4d, 16'h2c4e, 16'h2c4f, 16'h2c50, 16'h2c51, 16'h2c52, 16'h2c53, 16'h2c54, 16'h2c55, 16'h2c56, 16'h2c57, 16'h2c58, 16'h2c59, 16'h2c5a, 16'h2c5b, 16'h2c5c, 16'h2c5d, 16'h2c5e, 16'h2c5f, 16'h2c60, 16'h2c61, 16'h2c62, 16'h2c63, 16'h2c64, 16'h2c65, 16'h2c66, 16'h2c67, 16'h2c68, 16'h2c69, 16'h2c6a, 16'h2c6b, 16'h2c6c, 16'h2c6d, 16'h2c6e, 16'h2c6f, 16'h2c70, 16'h2c71, 16'h2c72, 16'h2c73},
                                {16'h2c74, 16'h2c75, 16'h2c76, 16'h2c77, 16'h2c78, 16'h2c79, 16'h2c7a, 16'h2c7b, 16'h2c7c, 16'h2c7d, 16'h2c7e, 16'h2c7f, 16'h2c80, 16'h2c81, 16'h2c82, 16'h2c83, 16'h2c84, 16'h2c85, 16'h2c86, 16'h2c87, 16'h2c88, 16'h2c89, 16'h2c8a, 16'h2c8b, 16'h2c8c, 16'h2c8d, 16'h2c8e, 16'h2c8f, 16'h2c90, 16'h2c91, 16'h2c92, 16'h2c93, 16'h2c94, 16'h2c95, 16'h2c96, 16'h2c97, 16'h2c98, 16'h2c99, 16'h2c9a, 16'h2c9b, 16'h2c9c, 16'h2c9d, 16'h2c9e, 16'h2c9f, 16'h2ca0, 16'h2ca1, 16'h2ca2, 16'h2ca3, 16'h2ca4, 16'h2ca5, 16'h2ca6, 16'h2ca7, 16'h2ca8, 16'h2ca9, 16'h2caa, 16'h2cab, 16'h2cac, 16'h2cad, 16'h2cae, 16'h2caf, 16'h2cb0, 16'h2cb1, 16'h2cb2, 16'h2cb3},
                                {16'h2cb4, 16'h2cb5, 16'h2cb6, 16'h2cb7, 16'h2cb8, 16'h2cb9, 16'h2cba, 16'h2cbb, 16'h2cbc, 16'h2cbd, 16'h2cbe, 16'h2cbf, 16'h2cc0, 16'h2cc1, 16'h2cc2, 16'h2cc3, 16'h2cc4, 16'h2cc5, 16'h2cc6, 16'h2cc7, 16'h2cc8, 16'h2cc9, 16'h2cca, 16'h2ccb, 16'h2ccc, 16'h2ccd, 16'h2cce, 16'h2ccf, 16'h2cd0, 16'h2cd1, 16'h2cd2, 16'h2cd3, 16'h2cd4, 16'h2cd5, 16'h2cd6, 16'h2cd7, 16'h2cd8, 16'h2cd9, 16'h2cda, 16'h2cdb, 16'h2cdc, 16'h2cdd, 16'h2cde, 16'h2cdf, 16'h2ce0, 16'h2ce1, 16'h2ce2, 16'h2ce3, 16'h2ce4, 16'h2ce5, 16'h2ce6, 16'h2ce7, 16'h2ce8, 16'h2ce9, 16'h2cea, 16'h2ceb, 16'h2cec, 16'h2ced, 16'h2cee, 16'h2cef, 16'h2cf0, 16'h2cf1, 16'h2cf2, 16'h2cf3},
                                {16'h2cf4, 16'h2cf5, 16'h2cf6, 16'h2cf7, 16'h2cf8, 16'h2cf9, 16'h2cfa, 16'h2cfb, 16'h2cfc, 16'h2cfd, 16'h2cfe, 16'h2cff, 16'h2d00, 16'h2d01, 16'h2d02, 16'h2d03, 16'h2d04, 16'h2d05, 16'h2d06, 16'h2d07, 16'h2d08, 16'h2d09, 16'h2d0a, 16'h2d0b, 16'h2d0c, 16'h2d0d, 16'h2d0e, 16'h2d0f, 16'h2d10, 16'h2d11, 16'h2d12, 16'h2d13, 16'h2d14, 16'h2d15, 16'h2d16, 16'h2d17, 16'h2d18, 16'h2d19, 16'h2d1a, 16'h2d1b, 16'h2d1c, 16'h2d1d, 16'h2d1e, 16'h2d1f, 16'h2d20, 16'h2d21, 16'h2d22, 16'h2d23, 16'h2d24, 16'h2d25, 16'h2d26, 16'h2d27, 16'h2d28, 16'h2d29, 16'h2d2a, 16'h2d2b, 16'h2d2c, 16'h2d2d, 16'h2d2e, 16'h2d2f, 16'h2d30, 16'h2d31, 16'h2d32, 16'h2d33},
                                {16'h2d34, 16'h2d35, 16'h2d36, 16'h2d37, 16'h2d38, 16'h2d39, 16'h2d3a, 16'h2d3b, 16'h2d3c, 16'h2d3d, 16'h2d3e, 16'h2d3f, 16'h2d40, 16'h2d41, 16'h2d42, 16'h2d43, 16'h2d44, 16'h2d45, 16'h2d46, 16'h2d47, 16'h2d48, 16'h2d49, 16'h2d4a, 16'h2d4b, 16'h2d4c, 16'h2d4d, 16'h2d4e, 16'h2d4f, 16'h2d50, 16'h2d51, 16'h2d52, 16'h2d53, 16'h2d54, 16'h2d55, 16'h2d56, 16'h2d57, 16'h2d58, 16'h2d59, 16'h2d5a, 16'h2d5b, 16'h2d5c, 16'h2d5d, 16'h2d5e, 16'h2d5f, 16'h2d60, 16'h2d61, 16'h2d62, 16'h2d63, 16'h2d64, 16'h2d65, 16'h2d66, 16'h2d67, 16'h2d68, 16'h2d69, 16'h2d6a, 16'h2d6b, 16'h2d6c, 16'h2d6d, 16'h2d6e, 16'h2d6f, 16'h2d70, 16'h2d71, 16'h2d72, 16'h2d73},
                                {16'h2d74, 16'h2d75, 16'h2d76, 16'h2d77, 16'h2d78, 16'h2d79, 16'h2d7a, 16'h2d7b, 16'h2d7c, 16'h2d7d, 16'h2d7e, 16'h2d7f, 16'h2d80, 16'h2d81, 16'h2d82, 16'h2d83, 16'h2d84, 16'h2d85, 16'h2d86, 16'h2d87, 16'h2d88, 16'h2d89, 16'h2d8a, 16'h2d8b, 16'h2d8c, 16'h2d8d, 16'h2d8e, 16'h2d8f, 16'h2d90, 16'h2d91, 16'h2d92, 16'h2d93, 16'h2d94, 16'h2d95, 16'h2d96, 16'h2d97, 16'h2d98, 16'h2d99, 16'h2d9a, 16'h2d9b, 16'h2d9c, 16'h2d9d, 16'h2d9e, 16'h2d9f, 16'h2da0, 16'h2da1, 16'h2da2, 16'h2da3, 16'h2da4, 16'h2da5, 16'h2da6, 16'h2da7, 16'h2da8, 16'h2da9, 16'h2daa, 16'h2dab, 16'h2dac, 16'h2dad, 16'h2dae, 16'h2daf, 16'h2db0, 16'h2db1, 16'h2db2, 16'h2db3},
                                {16'h2db4, 16'h2db5, 16'h2db6, 16'h2db7, 16'h2db8, 16'h2db9, 16'h2dba, 16'h2dbb, 16'h2dbc, 16'h2dbd, 16'h2dbe, 16'h2dbf, 16'h2dc0, 16'h2dc1, 16'h2dc2, 16'h2dc3, 16'h2dc4, 16'h2dc5, 16'h2dc6, 16'h2dc7, 16'h2dc8, 16'h2dc9, 16'h2dca, 16'h2dcb, 16'h2dcc, 16'h2dcd, 16'h2dce, 16'h2dcf, 16'h2dd0, 16'h2dd1, 16'h2dd2, 16'h2dd3, 16'h2dd4, 16'h2dd5, 16'h2dd6, 16'h2dd7, 16'h2dd8, 16'h2dd9, 16'h2dda, 16'h2ddb, 16'h2ddc, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd},
                                {16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd},
                                {16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd},
                                {16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd},
                                {16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd},
                                {16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd},
                                {16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd},
                                {16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd},
                                {16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd},
                                {16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd},
                                {16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd},
                                {16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd},
                                {16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd},
                                {16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd},
                                {16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd},
                                {16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd},
                                {16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd},
                                {16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd},
                                {16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd},
                                {16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd},
                                {16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd},
                                {16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd},
                                {16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd},
                                {16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd},
                                {16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd},
                                {16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd},
                                {16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd},
                                {16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddd, 16'h2ddc, 16'h2ddb, 16'h2dda, 16'h2dd9, 16'h2dd8, 16'h2dd7, 16'h2dd6, 16'h2dd5, 16'h2dd4, 16'h2dd3, 16'h2dd2, 16'h2dd1, 16'h2dd0, 16'h2dcf, 16'h2dce, 16'h2dcd, 16'h2dcc, 16'h2dcb, 16'h2dca, 16'h2dc9, 16'h2dc8, 16'h2dc7, 16'h2dc6, 16'h2dc5, 16'h2dc4, 16'h2dc3, 16'h2dc2, 16'h2dc1, 16'h2dc0, 16'h2dbf, 16'h2dbe, 16'h2dbd, 16'h2dbc, 16'h2dbb, 16'h2dba, 16'h2db9, 16'h2db8, 16'h2db7, 16'h2db6, 16'h2db5, 16'h2db4, 16'h2db3, 16'h2db2, 16'h2db1},
                                {16'h2db0, 16'h2daf, 16'h2dae, 16'h2dad, 16'h2dac, 16'h2dab, 16'h2daa, 16'h2da9, 16'h2da8, 16'h2da7, 16'h2da6, 16'h2da5, 16'h2da4, 16'h2da3, 16'h2da2, 16'h2da1, 16'h2da0, 16'h2d9f, 16'h2d9e, 16'h2d9d, 16'h2d9c, 16'h2d9b, 16'h2d9a, 16'h2d99, 16'h2d98, 16'h2d97, 16'h2d96, 16'h2d95, 16'h2d94, 16'h2d93, 16'h2d92, 16'h2d91, 16'h2d90, 16'h2d8f, 16'h2d8e, 16'h2d8d, 16'h2d8c, 16'h2d8b, 16'h2d8a, 16'h2d89, 16'h2d88, 16'h2d87, 16'h2d86, 16'h2d85, 16'h2d84, 16'h2d83, 16'h2d82, 16'h2d81, 16'h2d80, 16'h2d7f, 16'h2d7e, 16'h2d7d, 16'h2d7c, 16'h2d7b, 16'h2d7a, 16'h2d79, 16'h2d78, 16'h2d77, 16'h2d76, 16'h2d75, 16'h2d74, 16'h2d73, 16'h2d72, 16'h2d71},
                                {16'h2d70, 16'h2d6f, 16'h2d6e, 16'h2d6d, 16'h2d6c, 16'h2d6b, 16'h2d6a, 16'h2d69, 16'h2d68, 16'h2d67, 16'h2d66, 16'h2d65, 16'h2d64, 16'h2d63, 16'h2d62, 16'h2d61, 16'h2d60, 16'h2d5f, 16'h2d5e, 16'h2d5d, 16'h2d5c, 16'h2d5b, 16'h2d5a, 16'h2d59, 16'h2d58, 16'h2d57, 16'h2d56, 16'h2d55, 16'h2d54, 16'h2d53, 16'h2d52, 16'h2d51, 16'h2d50, 16'h2d4f, 16'h2d4e, 16'h2d4d, 16'h2d4c, 16'h2d4b, 16'h2d4a, 16'h2d49, 16'h2d48, 16'h2d47, 16'h2d46, 16'h2d45, 16'h2d44, 16'h2d43, 16'h2d42, 16'h2d41, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40},
                                {16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40},
                                {16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40},
                                {16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40},
                                {16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40},
                                {16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40},
                                {16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40},
                                {16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40},
                                {16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40},
                                {16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40},
                                {16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40},
                                {16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40},
                                {16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40},
                                {16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40},
                                {16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40},
                                {16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40},
                                {16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40},
                                {16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40},
                                {16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40},
                                {16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40},
                                {16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40},
                                {16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40},
                                {16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40},
                                {16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40},
                                {16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40},
                                {16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40},
                                {16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40},
                                {16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d40, 16'h2d3f, 16'h2d3e, 16'h2d3d, 16'h2d3c, 16'h2d3b, 16'h2d3a, 16'h2d39, 16'h2d38, 16'h2d37, 16'h2d36, 16'h2d35, 16'h2d34, 16'h2d33, 16'h2d32, 16'h2d31, 16'h2d30, 16'h2d2f, 16'h2d2e, 16'h2d2d, 16'h2d2c, 16'h2d2b, 16'h2d2a, 16'h2d29, 16'h2d28, 16'h2d27, 16'h2d26, 16'h2d25, 16'h2d24, 16'h2d23, 16'h2d22, 16'h2d21, 16'h2d20, 16'h2d1f, 16'h2d1e, 16'h2d1d, 16'h2d1c, 16'h2d1b, 16'h2d1a, 16'h2d19},
                                {16'h2d18, 16'h2d17, 16'h2d16, 16'h2d15, 16'h2d14, 16'h2d13, 16'h2d12, 16'h2d11, 16'h2d10, 16'h2d0f, 16'h2d0e, 16'h2d0d, 16'h2d0c, 16'h2d0b, 16'h2d0a, 16'h2d09, 16'h2d08, 16'h2d07, 16'h2d06, 16'h2d05, 16'h2d04, 16'h2d03, 16'h2d02, 16'h2d01, 16'h2d00, 16'h2cff, 16'h2cfe, 16'h2cfd, 16'h2cfc, 16'h2cfb, 16'h2cfa, 16'h2cf9, 16'h2cf8, 16'h2cf7, 16'h2cf6, 16'h2cf5, 16'h2cf4, 16'h2cf3, 16'h2cf2, 16'h2cf1, 16'h2cf0, 16'h2cef, 16'h2cee, 16'h2ced, 16'h2cec, 16'h2ceb, 16'h2cea, 16'h2ce9, 16'h2ce8, 16'h2ce7, 16'h2ce6, 16'h2ce5, 16'h2ce4, 16'h2ce3, 16'h2ce2, 16'h2ce1, 16'h2ce0, 16'h2cdf, 16'h2cde, 16'h2cdd, 16'h2cdc, 16'h2cdb, 16'h2cda, 16'h2cd9},
                                {16'h2cd8, 16'h2cd7, 16'h2cd6, 16'h2cd5, 16'h2cd4, 16'h2cd3, 16'h2cd2, 16'h2cd1, 16'h2cd0, 16'h2ccf, 16'h2cce, 16'h2ccd, 16'h2ccc, 16'h2ccb, 16'h2cca, 16'h2cc9, 16'h2cc8, 16'h2cc7, 16'h2cc6, 16'h2cc5, 16'h2cc4, 16'h2cc3, 16'h2cc2, 16'h2cc1, 16'h2cc0, 16'h2cbf, 16'h2cbe, 16'h2cbd, 16'h2cbc, 16'h2cbb, 16'h2cba, 16'h2cb9, 16'h2cb8, 16'h2cb7, 16'h2cb6, 16'h2cb5, 16'h2cb4, 16'h2cb3, 16'h2cb2, 16'h2cb1, 16'h2cb0, 16'h2caf, 16'h2cae, 16'h2cad, 16'h2cac, 16'h2cab, 16'h2caa, 16'h2ca9, 16'h2ca8, 16'h2ca7, 16'h2ca6, 16'h2ca5, 16'h2ca4, 16'h2ca3, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2},
                                {16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2},
                                {16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2},
                                {16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2},
                                {16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2},
                                {16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2},
                                {16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2},
                                {16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2},
                                {16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2},
                                {16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2},
                                {16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2},
                                {16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2},
                                {16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2},
                                {16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2},
                                {16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2},
                                {16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2},
                                {16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2},
                                {16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2},
                                {16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2},
                                {16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2},
                                {16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2},
                                {16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2},
                                {16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca2, 16'h2ca1, 16'h2ca0, 16'h2c9f, 16'h2c9e, 16'h2c9d, 16'h2c9c, 16'h2c9b, 16'h2c9a, 16'h2c99, 16'h2c98, 16'h2c97, 16'h2c96, 16'h2c95, 16'h2c94, 16'h2c93, 16'h2c92, 16'h2c91, 16'h2c90, 16'h2c8f, 16'h2c8e, 16'h2c8d, 16'h2c8c, 16'h2c8b, 16'h2c8a, 16'h2c89, 16'h2c88, 16'h2c87, 16'h2c86, 16'h2c85, 16'h2c84, 16'h2c83, 16'h2c82, 16'h2c81, 16'h2c80, 16'h2c7f, 16'h2c7e, 16'h2c7d, 16'h2c7c, 16'h2c7b, 16'h2c7a, 16'h2c79, 16'h2c78, 16'h2c77, 16'h2c76, 16'h2c75, 16'h2c74, 16'h2c73, 16'h2c72, 16'h2c71, 16'h2c70, 16'h2c6f, 16'h2c6e, 16'h2c6d, 16'h2c6c, 16'h2c6b, 16'h2c6a, 16'h2c69, 16'h2c68},
                                {16'h2c67, 16'h2c66, 16'h2c65, 16'h2c64, 16'h2c63, 16'h2c62, 16'h2c61, 16'h2c60, 16'h2c5f, 16'h2c5e, 16'h2c5d, 16'h2c5c, 16'h2c5b, 16'h2c5a, 16'h2c59, 16'h2c58, 16'h2c57, 16'h2c56, 16'h2c55, 16'h2c54, 16'h2c53, 16'h2c52, 16'h2c51, 16'h2c50, 16'h2c4f, 16'h2c4e, 16'h2c4d, 16'h2c4c, 16'h2c4b, 16'h2c4a, 16'h2c49, 16'h2c48, 16'h2c47, 16'h2c46, 16'h2c45, 16'h2c44, 16'h2c43, 16'h2c42, 16'h2c41, 16'h2c40, 16'h2c3f, 16'h2c3e, 16'h2c3d, 16'h2c3c, 16'h2c3b, 16'h2c3a, 16'h2c39, 16'h2c38, 16'h2c37, 16'h2c36, 16'h2c35, 16'h2c34, 16'h2c33, 16'h2c32, 16'h2c31, 16'h2c30, 16'h2c2f, 16'h2c2e, 16'h2c2d, 16'h2c2c, 16'h2c2b, 16'h2c2a, 16'h2c29, 16'h2c28},
                                {16'h2c27, 16'h2c26, 16'h2c25, 16'h2c24, 16'h2c23, 16'h2c22, 16'h2c21, 16'h2c20, 16'h2c1f, 16'h2c1e, 16'h2c1d, 16'h2c1c, 16'h2c1b, 16'h2c1a, 16'h2c19, 16'h2c18, 16'h2c17, 16'h2c16, 16'h2c15, 16'h2c14, 16'h2c13, 16'h2c12, 16'h2c11, 16'h2c10, 16'h2c0f, 16'h2c0e, 16'h2c0d, 16'h2c0c, 16'h2c0b, 16'h2c0a, 16'h2c09, 16'h2c08, 16'h2c07, 16'h2c06, 16'h2c05, 16'h2c04, 16'h2c03, 16'h2c02, 16'h2c01, 16'h2c00, 16'h2bff, 16'h2bfe, 16'h2bfd, 16'h2bfc, 16'h2bfb, 16'h2bfa, 16'h2bf9, 16'h2bf8, 16'h2bf7, 16'h2bf6, 16'h2bf5, 16'h2bf4, 16'h2bf3, 16'h2bf2, 16'h2bf1, 16'h2bf0, 16'h2bef, 16'h2bee, 16'h2bed, 16'h2bec, 16'h2beb, 16'h2bea, 16'h2be9, 16'h2be8},
                                {16'h2be7, 16'h2be6, 16'h2be5, 16'h2be4, 16'h2be3, 16'h2be2, 16'h2be1, 16'h2be0, 16'h2bdf, 16'h2bde, 16'h2bdd, 16'h2bdc, 16'h2bdb, 16'h2bda, 16'h2bd9, 16'h2bd8, 16'h2bd7, 16'h2bd6, 16'h2bd5, 16'h2bd4, 16'h2bd3, 16'h2bd2, 16'h2bd1, 16'h2bd0, 16'h2bcf, 16'h2bce, 16'h2bcd, 16'h2bcc, 16'h2bcb, 16'h2bca, 16'h2bc9, 16'h2bc8, 16'h2bc7, 16'h2bc6, 16'h2bc5, 16'h2bc4, 16'h2bc3, 16'h2bc2, 16'h2bc1, 16'h2bc0, 16'h2bbf, 16'h2bbe, 16'h2bbd, 16'h2bbc, 16'h2bbb, 16'h2bba, 16'h2bb9, 16'h2bb8, 16'h2bb7, 16'h2bb6, 16'h2bb5, 16'h2bb4, 16'h2bb3, 16'h2bb2, 16'h2bb1, 16'h2bb0, 16'h2baf, 16'h2bae, 16'h2bad, 16'h2bac, 16'h2bab, 16'h2baa, 16'h2ba9, 16'h2ba8},
                                {16'h2ba7, 16'h2ba6, 16'h2ba5, 16'h2ba4, 16'h2ba3, 16'h2ba2, 16'h2ba1, 16'h2ba0, 16'h2b9f, 16'h2b9e, 16'h2b9d, 16'h2b9c, 16'h2b9b, 16'h2b9a, 16'h2b99, 16'h2b98, 16'h2b97, 16'h2b96, 16'h2b95, 16'h2b94, 16'h2b93, 16'h2b92, 16'h2b91, 16'h2b90, 16'h2b8f, 16'h2b8e, 16'h2b8d, 16'h2b8c, 16'h2b8b, 16'h2b8a, 16'h2b89, 16'h2b88, 16'h2b87, 16'h2b86, 16'h2b85, 16'h2b84, 16'h2b83, 16'h2b82, 16'h2b81, 16'h2b80, 16'h2b7f, 16'h2b7e, 16'h2b7d, 16'h2b7c, 16'h2b7b, 16'h2b7a, 16'h2b79, 16'h2b78, 16'h2b77, 16'h2b76, 16'h2b75, 16'h2b74, 16'h2b73, 16'h2b72, 16'h2b71, 16'h2b70, 16'h2b6f, 16'h2b6e, 16'h2b6d, 16'h2b6c, 16'h2b6b, 16'h2b6a, 16'h2b69, 16'h2b68},
                                {16'h2b67, 16'h2b66, 16'h2b65, 16'h2b64, 16'h2b63, 16'h2b62, 16'h2b61, 16'h2b60, 16'h2b5f, 16'h2b5e, 16'h2b5d, 16'h2b5c, 16'h2b5b, 16'h2b5a, 16'h2b59, 16'h2b58, 16'h2b57, 16'h2b56, 16'h2b55, 16'h2b54, 16'h2b71, 16'h2b72, 16'h2b73, 16'h2b74, 16'h2b75, 16'h2b76, 16'h2b77, 16'h2b78, 16'h2b79, 16'h2b7a, 16'h2b7b, 16'h2b7c, 16'h2b7d, 16'h2b7e, 16'h2b7f, 16'h2b80, 16'h2b81, 16'h2b82, 16'h2b83, 16'h2b84, 16'h2b85, 16'h2b86, 16'h2b87, 16'h2b88, 16'h2b89, 16'h2b8a, 16'h2b8b, 16'h2b8c, 16'h2b8d, 16'h2b8e, 16'h2b8f, 16'h2b90, 16'h2b91, 16'h2b92, 16'h2b93, 16'h2b94, 16'h2b95, 16'h2b96, 16'h2b97, 16'h2b98, 16'h2b99, 16'h2b9a, 16'h2b9b, 16'h2b9c},
                                {16'h2b9d, 16'h2b9e, 16'h2b9f, 16'h2ba0, 16'h2ba1, 16'h2ba2, 16'h2ba3, 16'h2ba4, 16'h2ba5, 16'h2ba6, 16'h2ba7, 16'h2ba8, 16'h2ba9, 16'h2baa, 16'h2bab, 16'h2bac, 16'h2bad, 16'h2bae, 16'h2baf, 16'h2bb0, 16'h2bb1, 16'h2bb2, 16'h2bb3, 16'h2bb4, 16'h2bb5, 16'h2bb6, 16'h2bb7, 16'h2bb8, 16'h2bb9, 16'h2bba, 16'h2bbb, 16'h2bbc, 16'h2bbd, 16'h2bbe, 16'h2bbf, 16'h2bc0, 16'h2bc1, 16'h2bc2, 16'h2bc3, 16'h2bc4, 16'h2bc5, 16'h2bc6, 16'h2bc7, 16'h2bc8, 16'h2bc9, 16'h2bca, 16'h2bcb, 16'h2bcc, 16'h2bcd, 16'h2bce, 16'h2bcf, 16'h2bd0, 16'h2bd1, 16'h2bd2, 16'h2bd3, 16'h2bd4, 16'h2bd5, 16'h2bd6, 16'h2bd7, 16'h2bd8, 16'h2bd9, 16'h2bda, 16'h2bdb, 16'h2bdc},
                                {16'h2bdd, 16'h2bde, 16'h2bdf, 16'h2be0, 16'h2be1, 16'h2be2, 16'h2be3, 16'h2be4, 16'h2be5, 16'h2be6, 16'h2be7, 16'h2be8, 16'h2be9, 16'h2bea, 16'h2beb, 16'h2bec, 16'h2bed, 16'h2bee, 16'h2bef, 16'h2bf0, 16'h2bf1, 16'h2bf2, 16'h2bf3, 16'h2bf4, 16'h2bf5, 16'h2bf6, 16'h2bf7, 16'h2bf8, 16'h2bf9, 16'h2bfa, 16'h2bfb, 16'h2bfc, 16'h2bfd, 16'h2bfe, 16'h2bff, 16'h2c00, 16'h2c01, 16'h2c02, 16'h2c03, 16'h2c04, 16'h2c05, 16'h2c06, 16'h2c07, 16'h2c08, 16'h2c09, 16'h2c0a, 16'h2c0b, 16'h2c0c, 16'h2c0d, 16'h2c0e, 16'h2c0f, 16'h2c10, 16'h2c11, 16'h2c12, 16'h2c13, 16'h2c14, 16'h2c15, 16'h2c16, 16'h2c17, 16'h2c18, 16'h2c19, 16'h2ac5, 16'h296c, 16'h2813},
                                {16'h26ba, 16'h2561, 16'h2408, 16'h22af, 16'h2156, 16'h1ffd, 16'h1ea4, 16'h1d4b, 16'h1bf2, 16'h1a99, 16'h1940, 16'h17e7, 16'h168e, 16'h1535, 16'h13dc, 16'h1283, 16'h126c, 16'h1248, 16'h1224, 16'h1200, 16'h11dc, 16'h11b8, 16'h1194, 16'h1170, 16'h114c, 16'h1128, 16'h1104, 16'h10e0, 16'h10bc, 16'h1098, 16'h1074, 16'h1050, 16'h102c, 16'h1008, 16'h0fe4, 16'h0fc0, 16'h0f9c, 16'h0f78, 16'h0f54, 16'h0f30, 16'h0f0c, 16'h0ee8, 16'h0ec4, 16'h0ea0, 16'h0e7c, 16'h0e58, 16'h0e34, 16'h0e10, 16'h0dec, 16'h0dc8, 16'h0da4, 16'h0d80, 16'h0d5c, 16'h0d38, 16'h0d14, 16'h0cf0, 16'h0ccc, 16'h0ca8, 16'h0c84, 16'h0c60, 16'h0c3c, 16'h0c18, 16'h0bf4, 16'h0bd0},
                                {16'h0bac, 16'h0b88, 16'h0b64, 16'h0b40, 16'h0b1c, 16'h0af8, 16'h0ad4, 16'h0ab0, 16'h0a8c, 16'h0a68, 16'h0a44, 16'h0a20, 16'h09fc, 16'h09d8, 16'h09b4, 16'h0990, 16'h096c, 16'h0948, 16'h0924, 16'h0900, 16'h08dc, 16'h08b8, 16'h0894, 16'h0870, 16'h084c, 16'h0828, 16'h0804, 16'h07e0, 16'h07bc, 16'h0798, 16'h0774, 16'h0750, 16'h072c, 16'h0708, 16'h06e4, 16'h06c0, 16'h069c, 16'h0678, 16'h0654, 16'h0630, 16'h060c, 16'h05e8, 16'h05c4, 16'h05a0, 16'h057c, 16'h0558, 16'h0534, 16'h0510, 16'h04ec, 16'h04c8, 16'h04a4, 16'h0480, 16'h045c, 16'h0438, 16'h0414, 16'h03f0, 16'h03cc, 16'h03a8, 16'h0384, 16'h0360, 16'h033c, 16'h0318, 16'h02f4, 16'h02d0},
                                {16'h02ac, 16'h0288, 16'h0264, 16'h0240, 16'h021c, 16'h01f8, 16'h01d4, 16'h01b0, 16'h018c, 16'h0168, 16'h0144, 16'h0120, 16'h00fc, 16'h00d8, 16'h00b4, 16'h0090, 16'h006c, 16'h0048, 16'h0024, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000},
                                {16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000},
                                {16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000},
                                {16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000},
                                {16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000},
                                {16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000},
                                {16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000},
                                {16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000},
                                {16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000},
                                {16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000},
                                {16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000},
                                {16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000},
                                {16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000},
                                {16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000},
                                {16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000},
                                {16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000},
                                {16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000},
                                {16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000},
                                {16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000},
                                {16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000},
                                {16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000},
                                {16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000},
                                {16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000},
                                {16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000},
                                {16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000},
                                {16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0001, 16'h0002, 16'h0003, 16'h0004, 16'h0005, 16'h0006, 16'h0007, 16'h0008, 16'h0009, 16'h000a, 16'h000b, 16'h000c, 16'h000d, 16'h000e, 16'h000f, 16'h0010, 16'h0011, 16'h0012, 16'h0013, 16'h0014, 16'h0015, 16'h0016, 16'h0017, 16'h0018, 16'h0019, 16'h001a, 16'h001b, 16'h001c, 16'h001d, 16'h001e, 16'h001f, 16'h0020, 16'h0021, 16'h0022, 16'h0023, 16'h0024, 16'h0025, 16'h0026, 16'h0027, 16'h0028, 16'h0029, 16'h002a, 16'h002b, 16'h002c, 16'h002d, 16'h002e, 16'h002f, 16'h0030, 16'h0031, 16'h0032},
                                {16'h0033, 16'h0034, 16'h0035, 16'h0036, 16'h0037, 16'h0038, 16'h0039, 16'h003a, 16'h003b, 16'h003c, 16'h003d, 16'h003e, 16'h003f, 16'h0040, 16'h0041, 16'h0042, 16'h0043, 16'h0044, 16'h0045, 16'h0046, 16'h0047, 16'h0048, 16'h0049, 16'h004a, 16'h004b, 16'h004c, 16'h004d, 16'h004e, 16'h004f, 16'h0050, 16'h0051, 16'h0052, 16'h0053, 16'h0054, 16'h0055, 16'h0056, 16'h0057, 16'h0058, 16'h0059, 16'h005a, 16'h005b, 16'h005c, 16'h005d, 16'h005e, 16'h005f, 16'h0060, 16'h0061, 16'h0062, 16'h0063, 16'h0064, 16'h0065, 16'h0066, 16'h0067, 16'h0068, 16'h0069, 16'h006a, 16'h006b, 16'h006c, 16'h006d, 16'h006e, 16'h006f, 16'h0070, 16'h0071, 16'h0072},
                                {16'h0073, 16'h0074, 16'h0075, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076},
                                {16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076},
                                {16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076},
                                {16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076},
                                {16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076},
                                {16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076},
                                {16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076},
                                {16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076},
                                {16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076},
                                {16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076},
                                {16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076},
                                {16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076},
                                {16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076},
                                {16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076},
                                {16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076},
                                {16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076},
                                {16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076},
                                {16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076},
                                {16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076},
                                {16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076},
                                {16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076},
                                {16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076},
                                {16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076},
                                {16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076},
                                {16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0077, 16'h0078},
                                {16'h0079, 16'h007a, 16'h007b, 16'h007c, 16'h007d, 16'h007e, 16'h007f, 16'h0080, 16'h0081, 16'h0082, 16'h0083, 16'h0084, 16'h0085, 16'h0086, 16'h0087, 16'h0088, 16'h0089, 16'h008a, 16'h008b, 16'h008c, 16'h008d, 16'h008e, 16'h008f, 16'h0090, 16'h0091, 16'h0092, 16'h0093, 16'h0094, 16'h0095, 16'h0096, 16'h0097, 16'h0098, 16'h0099, 16'h009a, 16'h009b, 16'h009c, 16'h009d, 16'h009e, 16'h009f, 16'h00a0, 16'h00a1, 16'h00a2, 16'h00a3, 16'h00a4, 16'h00a5, 16'h00a6, 16'h00a7, 16'h00a8, 16'h00a9, 16'h00aa, 16'h00ab, 16'h00ac, 16'h00ad, 16'h00ae, 16'h00af, 16'h00b0, 16'h00b1, 16'h00b2, 16'h00b3, 16'h00b4, 16'h00b5, 16'h00b6, 16'h00b7, 16'h00b8},
                                {16'h00b9, 16'h00ba, 16'h00bb, 16'h00bc, 16'h00bd, 16'h00be, 16'h00bf, 16'h00c0, 16'h00c1, 16'h00c2, 16'h00c3, 16'h00c4, 16'h00c5, 16'h00c6, 16'h00c7, 16'h00c8, 16'h00c9, 16'h00ca, 16'h00cb, 16'h00cc, 16'h00cd, 16'h00ce, 16'h00cf, 16'h00d0, 16'h00d1, 16'h00d2, 16'h00d3, 16'h00d4, 16'h00d5, 16'h00d6, 16'h00d7, 16'h00d8, 16'h00d9, 16'h00da, 16'h00db, 16'h00dc, 16'h00dd, 16'h00de, 16'h00df, 16'h00e0, 16'h00e1, 16'h00e2, 16'h00e3, 16'h00e4, 16'h00e5, 16'h00e6, 16'h00e7, 16'h00e8, 16'h00e9, 16'h00ea, 16'h00eb, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec},
                                {16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec},
                                {16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec},
                                {16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec},
                                {16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec},
                                {16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec},
                                {16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec},
                                {16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec},
                                {16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec},
                                {16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec},
                                {16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec},
                                {16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec},
                                {16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec},
                                {16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec},
                                {16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec},
                                {16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec},
                                {16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec},
                                {16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec},
                                {16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec},
                                {16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec},
                                {16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec},
                                {16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec},
                                {16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec},
                                {16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec},
                                {16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec},
                                {16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ec, 16'h00ed, 16'h00ee, 16'h00ef, 16'h00f0, 16'h00f1, 16'h00f2, 16'h00f3, 16'h00f4, 16'h00f5, 16'h00f6, 16'h00f7, 16'h00f8, 16'h00f9, 16'h00fa, 16'h00fb, 16'h00fc, 16'h00fd},
                                {16'h00fe, 16'h00ff, 16'h0100, 16'h0101, 16'h0102, 16'h0103, 16'h0104, 16'h0105, 16'h0106, 16'h0107, 16'h0108, 16'h0109, 16'h010a, 16'h010b, 16'h010c, 16'h010d, 16'h010e, 16'h010f, 16'h0110, 16'h0111, 16'h0112, 16'h0113, 16'h0114, 16'h0115, 16'h0116, 16'h0117, 16'h0118, 16'h0119, 16'h011a, 16'h011b, 16'h011c, 16'h011d, 16'h011e, 16'h011f, 16'h0120, 16'h0121, 16'h0122, 16'h0123, 16'h0124, 16'h0125, 16'h0126, 16'h0127, 16'h0128, 16'h0129, 16'h012a, 16'h012b, 16'h012c, 16'h012d, 16'h012e, 16'h012f, 16'h0130, 16'h0131, 16'h0132, 16'h0133, 16'h0134, 16'h0135, 16'h0136, 16'h0137, 16'h0138, 16'h0139, 16'h013a, 16'h013b, 16'h013c, 16'h013d},
                                {16'h013e, 16'h013f, 16'h0140, 16'h0141, 16'h0142, 16'h0143, 16'h0144, 16'h0145, 16'h0146, 16'h0147, 16'h0148, 16'h0149, 16'h014a, 16'h014b, 16'h014c, 16'h014d, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e},
                                {16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e},
                                {16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e},
                                {16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e},
                                {16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e},
                                {16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e},
                                {16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e},
                                {16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e},
                                {16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e},
                                {16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e},
                                {16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e},
                                {16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e},
                                {16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e},
                                {16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e},
                                {16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e},
                                {16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e},
                                {16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e},
                                {16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e},
                                {16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e},
                                {16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e},
                                {16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e},
                                {16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014e, 16'h014d, 16'h014c, 16'h014b, 16'h014a, 16'h0149, 16'h0148, 16'h0147, 16'h0146, 16'h0145, 16'h0144, 16'h0143, 16'h0142, 16'h0141, 16'h0140},
                                {16'h013f, 16'h013e, 16'h013d, 16'h013c, 16'h013b, 16'h013a, 16'h0139, 16'h0138, 16'h0137, 16'h0136, 16'h0135, 16'h0134, 16'h0133, 16'h0132, 16'h0131, 16'h0130, 16'h012f, 16'h012e, 16'h012d, 16'h012c, 16'h012b, 16'h012a, 16'h0129, 16'h0128, 16'h0127, 16'h0126, 16'h0125, 16'h0124, 16'h0123, 16'h0122, 16'h0121, 16'h0120, 16'h011f, 16'h011e, 16'h011d, 16'h011c, 16'h011b, 16'h011a, 16'h0119, 16'h0118, 16'h0117, 16'h0116, 16'h0115, 16'h0114, 16'h0113, 16'h0112, 16'h0111, 16'h0110, 16'h010f, 16'h010e, 16'h010d, 16'h010c, 16'h010b, 16'h010a, 16'h0109, 16'h0108, 16'h0107, 16'h0106, 16'h0105, 16'h0104, 16'h0103, 16'h0102, 16'h0101, 16'h0100},
                                {16'h00ff, 16'h00fe, 16'h00fd, 16'h00fc, 16'h00fb, 16'h00fa, 16'h00f9, 16'h00f8, 16'h00f7, 16'h00f6, 16'h00f5, 16'h00f4, 16'h00f3, 16'h00f2, 16'h00f1, 16'h00f0, 16'h00ef, 16'h00ee, 16'h00ed, 16'h00ec, 16'h00eb, 16'h00ea, 16'h00e9, 16'h00e8, 16'h00e7, 16'h00e6, 16'h00e5, 16'h00e4, 16'h00e3, 16'h00e2, 16'h00e1, 16'h00e0, 16'h00df, 16'h00de, 16'h00dd, 16'h00dc, 16'h00db, 16'h00da, 16'h00d9, 16'h00d8, 16'h00d7, 16'h00d6, 16'h00d5, 16'h00d4, 16'h00d3, 16'h00d2, 16'h00d1, 16'h00d0, 16'h00cf, 16'h00ce, 16'h00cd, 16'h00cc, 16'h00cb, 16'h00ca, 16'h00c9, 16'h00c8, 16'h00c7, 16'h00c6, 16'h00c5, 16'h00c4, 16'h00c3, 16'h00c2, 16'h00c1, 16'h00c0},
                                {16'h00bf, 16'h00be, 16'h00bd, 16'h00bc, 16'h00bb, 16'h00ba, 16'h00b9, 16'h00b8, 16'h00b7, 16'h00b6, 16'h00b5, 16'h00b4, 16'h00b3, 16'h00b2, 16'h00b1, 16'h00b0, 16'h00af, 16'h00ae, 16'h00ad, 16'h00ac, 16'h00ab, 16'h00aa, 16'h00a9, 16'h00a8, 16'h00a7, 16'h00a6, 16'h00a5, 16'h00a4, 16'h00a3, 16'h00a2, 16'h00a1, 16'h00a0, 16'h009f, 16'h009e, 16'h009d, 16'h009c, 16'h009b, 16'h009a, 16'h0099, 16'h0098, 16'h0097, 16'h0096, 16'h0095, 16'h0094, 16'h0093, 16'h0092, 16'h0091, 16'h0090, 16'h008f, 16'h008e, 16'h008d, 16'h008c, 16'h008b, 16'h008a, 16'h0089, 16'h0088, 16'h0087, 16'h0086, 16'h0085, 16'h0084, 16'h0083, 16'h0082, 16'h0081, 16'h0080},
                                {16'h007f, 16'h007e, 16'h007d, 16'h007c, 16'h007b, 16'h007a, 16'h0079, 16'h0078, 16'h0077, 16'h0076, 16'h0075, 16'h0074, 16'h0073, 16'h0072, 16'h0071, 16'h0070, 16'h006f, 16'h006e, 16'h006d, 16'h006c, 16'h006b, 16'h006a, 16'h0069, 16'h0068, 16'h0067, 16'h0066, 16'h0065, 16'h0064, 16'h0063, 16'h0062, 16'h0061, 16'h0060, 16'h005f, 16'h005e, 16'h005d, 16'h005c, 16'h005b, 16'h005a, 16'h0059, 16'h0058, 16'h0057, 16'h0056, 16'h0055, 16'h0054, 16'h0053, 16'h0052, 16'h0051, 16'h0050, 16'h004f, 16'h004e, 16'h004d, 16'h004c, 16'h004b, 16'h004a, 16'h0049, 16'h0048, 16'h0047, 16'h0046, 16'h0045, 16'h0044, 16'h0043, 16'h0042, 16'h0041, 16'h0040},
                                {16'h003f, 16'h003e, 16'h003d, 16'h003c, 16'h003b, 16'h003a, 16'h0039, 16'h0038, 16'h0037, 16'h0036, 16'h0035, 16'h0034, 16'h0033, 16'h0032, 16'h0031, 16'h0030, 16'h002f, 16'h002e, 16'h002d, 16'h002c, 16'h002b, 16'h002a, 16'h0029, 16'h0028, 16'h0027, 16'h0026, 16'h0025, 16'h0024, 16'h0023, 16'h0022, 16'h0021, 16'h0020, 16'h001f, 16'h001e, 16'h001d, 16'h001c, 16'h001b, 16'h001a, 16'h0019, 16'h0018, 16'h0017, 16'h0016, 16'h0015, 16'h0014, 16'h0013, 16'h0012, 16'h0011, 16'h0010, 16'h000f, 16'h000e, 16'h000d, 16'h000c, 16'h000b, 16'h000a, 16'h0009, 16'h0008, 16'h0007, 16'h0006, 16'h0005, 16'h0004, 16'h0003, 16'h0002, 16'h0001, 16'h0000}};
    DAC_Interface DUT (.clk(clk), .rst(rst),
                       .fresh_bits(fresh_bits),
                       .halt(1'b0),
                       .dac0_rdy(dac0_rdy),
                       .dac_batch(dac_batch),
                       .valid_dac_batch(valid_dac_batch),
                       .valid_dac_edge(valid_dac_edge),
                       .pwl_dma_if(pwl_dma_if));

    edetect #(.DATA_WIDTH(32))
    correct_ed(.clk(clk), .rst(rst),
               .val(correct_vals),
               .comb_posedge_out(correct_edge));
    always_comb begin
        for (int i = 0; i < `BATCH_SAMPLES; i++) begin
            dac_samples[i] = dac_batch[`SAMPLE_WIDTH*i+:`SAMPLE_WIDTH];
        end 
    end
    logic[31:0] test1, test2;
    assign test1 = `MAPPED_ID_CEILING;
    assign test2 = `MEM_SIZE-`MAPPED_ID_CEILING;
    always_ff@(posedge clk) begin
        if (rst) begin 
            {fresh_bits, pwl_dma_if.last, pwl_dma_if.data, pwl_dma_if.valid} <= 0;
            {exp_i,correct_vals} <= 0;
            timer <= 100;
            testState <= SEND;
        end
        else begin
            case(testState)
                SEND: begin 
                    if (timer == 100) fresh_bits[`PWL_PREP_ID] <= 1;
                    if (timer == 50) timer <= 0;
                    if (timer > 50) timer <= timer - 1;
                    else begin
                        if (timer == 0) begin 
                            timer <= 1; 
                            pwl_dma_if.valid <= 1; 
                            pwl_dma_if.data = dma_buff[0];
                            pwl_dma_if.last <= 0; 
                        end 
                        else if (timer < NUM_OF_POINTS) begin
                            if (pwl_dma_if.ready) begin
                                pwl_dma_if.data = dma_buff[timer];
                                if (timer == NUM_OF_POINTS-1) pwl_dma_if.last <= 1; 
                                timer <= timer + 1;
                            end 
                        end
                        else if (timer == NUM_OF_POINTS && pwl_dma_if.ready) begin
                            {pwl_dma_if.last, pwl_dma_if.data, pwl_dma_if.valid} <= 0;
                            timer <= 0; 
                            testState <= CHECK;
                        end
                    end
                end 
                CHECK: begin
                    if (exp_i == DUT.pwl_gen.wave_lines_stored) begin
                        exp_i <= 0; 
                        testState <= IDLE; 
                    end else begin
                        if (valid_dac_batch) begin
                            exp_i <= exp_i + 1;
                            if (curr_expected_batch == dac_samples) correct_vals <= correct_vals + 1; 
                            else correct_vals <= correct_vals - 1; 
                        end
                    end 
                end 
            endcase 

            if (fresh_bits) begin
                if (DUT.state_rdy) fresh_bits <= 0; 
            end 

            if (correct_edge == 1) begin 
                $write("%c[1;32m",27); 
                $write("t%0d+ ",exp_i);
                $write("%c[0m",27); 
            end else 
            if (correct_edge == 2) begin 
                $write("%c[1;31m",27); 
                $write("t%0d- ",exp_i);
                $write("%c[0m",27); 
            end 
        end
    end
    

    always begin
        #5;  
        clk = !clk;
    end

    initial begin
        $dumpfile("pwl2_tb.vcd");
        $dumpvars(0,pwl2_tb); 
        clk = 1;
        rst = 0;
        `flash_sig(rst); 
        #1000;
        while (testState != IDLE) #10;
        #70000;
        $finish;
    end 

endmodule 

`default_nettype wire
