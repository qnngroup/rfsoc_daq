// segmented_buffer_tb.sv - Reed Foster
// Tasks and driver submodules to verify segmented buffer


`timescale 1ns/1ps
module segmented_buffer_tb #(
  parameter int DISC_MAX_DELAY_CYCLES,
  parameter int BUFFER_READ_LATENCY
) (
);
endmodule


